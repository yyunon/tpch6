-- Copyright 2018-2019 Delft University of Technology
--
-- Licensed under the Apache License, Version 2.0 (the "License");
-- you may not use this file except in compliance with the License.
-- You may obtain a copy of the License at
--
--     http://www.apache.org/licenses/LICENSE-2.0
--
-- Unless required by applicable law or agreed to in writing, software
-- distributed under the License is distributed on an "AS IS" BASIS,
-- WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
-- See the License for the specific language governing permissions and
-- limitations under the License.
--
-- This file was generated by Fletchgen. Modify this file at your own risk.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.Interconnect_pkg.all;

entity Forecast_Mantle is
  generic (
    INDEX_WIDTH        : integer := 32;
    TAG_WIDTH          : integer := 1;
    BUS_ADDR_WIDTH     : integer := 64;
    BUS_DATA_WIDTH     : integer := 512;
    BUS_LEN_WIDTH      : integer := 8;
    BUS_BURST_STEP_LEN : integer := 1;
    BUS_BURST_MAX_LEN  : integer := 16
  );
  port (
    bcd_clk           : in  std_logic;
    bcd_reset         : in  std_logic;
    kcd_clk           : in  std_logic;
    kcd_reset         : in  std_logic;
    mmio_awvalid      : in  std_logic;
    mmio_awready      : out std_logic;
    mmio_awaddr       : in  std_logic_vector(31 downto 0);
    mmio_wvalid       : in  std_logic;
    mmio_wready       : out std_logic;
    mmio_wdata        : in  std_logic_vector(31 downto 0);
    mmio_wstrb        : in  std_logic_vector(3 downto 0);
    mmio_bvalid       : out std_logic;
    mmio_bready       : in  std_logic;
    mmio_bresp        : out std_logic_vector(1 downto 0);
    mmio_arvalid      : in  std_logic;
    mmio_arready      : out std_logic;
    mmio_araddr       : in  std_logic_vector(31 downto 0);
    mmio_rvalid       : out std_logic;
    mmio_rready       : in  std_logic;
    mmio_rdata        : out std_logic_vector(31 downto 0);
    mmio_rresp        : out std_logic_vector(1 downto 0);
    rd_mst_rreq_valid : out std_logic;
    rd_mst_rreq_ready : in  std_logic;
    rd_mst_rreq_addr  : out std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
    rd_mst_rreq_len   : out std_logic_vector(BUS_LEN_WIDTH-1 downto 0);
    rd_mst_rdat_valid : in  std_logic;
    rd_mst_rdat_ready : out std_logic;
    rd_mst_rdat_data  : in  std_logic_vector(BUS_DATA_WIDTH-1 downto 0);
    rd_mst_rdat_last  : in  std_logic
  );
end entity;

architecture Implementation of Forecast_Mantle is
  component Forecast_Nucleus is
    generic (
      INDEX_WIDTH                    : integer := 32;
      TAG_WIDTH                      : integer := 1;
      L_QUANTITY_BUS_ADDR_WIDTH      : integer := 64;
      L_EXTENDEDPRICE_BUS_ADDR_WIDTH : integer := 64;
      L_DISCOUNT_BUS_ADDR_WIDTH      : integer := 64;
      L_SHIPDATE_BUS_ADDR_WIDTH      : integer := 64
    );
    port (
      kcd_clk                      : in  std_logic;
      kcd_reset                    : in  std_logic;
      mmio_awvalid                 : in  std_logic;
      mmio_awready                 : out std_logic;
      mmio_awaddr                  : in  std_logic_vector(31 downto 0);
      mmio_wvalid                  : in  std_logic;
      mmio_wready                  : out std_logic;
      mmio_wdata                   : in  std_logic_vector(31 downto 0);
      mmio_wstrb                   : in  std_logic_vector(3 downto 0);
      mmio_bvalid                  : out std_logic;
      mmio_bready                  : in  std_logic;
      mmio_bresp                   : out std_logic_vector(1 downto 0);
      mmio_arvalid                 : in  std_logic;
      mmio_arready                 : out std_logic;
      mmio_araddr                  : in  std_logic_vector(31 downto 0);
      mmio_rvalid                  : out std_logic;
      mmio_rready                  : in  std_logic;
      mmio_rdata                   : out std_logic_vector(31 downto 0);
      mmio_rresp                   : out std_logic_vector(1 downto 0);
      l_quantity_valid             : in  std_logic;
      l_quantity_ready             : out std_logic;
      l_quantity_dvalid            : in  std_logic;
      l_quantity_last              : in  std_logic;
      l_quantity                   : in  std_logic_vector(63 downto 0);
      l_extendedprice_valid        : in  std_logic;
      l_extendedprice_ready        : out std_logic;
      l_extendedprice_dvalid       : in  std_logic;
      l_extendedprice_last         : in  std_logic;
      l_extendedprice              : in  std_logic_vector(63 downto 0);
      l_discount_valid             : in  std_logic;
      l_discount_ready             : out std_logic;
      l_discount_dvalid            : in  std_logic;
      l_discount_last              : in  std_logic;
      l_discount                   : in  std_logic_vector(63 downto 0);
      l_shipdate_valid             : in  std_logic;
      l_shipdate_ready             : out std_logic;
      l_shipdate_dvalid            : in  std_logic;
      l_shipdate_last              : in  std_logic;
      l_shipdate                   : in  std_logic_vector(63 downto 0);
      l_quantity_unl_valid         : in  std_logic;
      l_quantity_unl_ready         : out std_logic;
      l_quantity_unl_tag           : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      l_extendedprice_unl_valid    : in  std_logic;
      l_extendedprice_unl_ready    : out std_logic;
      l_extendedprice_unl_tag      : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      l_discount_unl_valid         : in  std_logic;
      l_discount_unl_ready         : out std_logic;
      l_discount_unl_tag           : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      l_shipdate_unl_valid         : in  std_logic;
      l_shipdate_unl_ready         : out std_logic;
      l_shipdate_unl_tag           : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      l_quantity_cmd_valid         : out std_logic;
      l_quantity_cmd_ready         : in  std_logic;
      l_quantity_cmd_firstIdx      : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      l_quantity_cmd_lastIdx       : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      l_quantity_cmd_ctrl          : out std_logic_vector(L_QUANTITY_BUS_ADDR_WIDTH-1 downto 0);
      l_quantity_cmd_tag           : out std_logic_vector(TAG_WIDTH-1 downto 0);
      l_extendedprice_cmd_valid    : out std_logic;
      l_extendedprice_cmd_ready    : in  std_logic;
      l_extendedprice_cmd_firstIdx : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      l_extendedprice_cmd_lastIdx  : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      l_extendedprice_cmd_ctrl     : out std_logic_vector(L_EXTENDEDPRICE_BUS_ADDR_WIDTH-1 downto 0);
      l_extendedprice_cmd_tag      : out std_logic_vector(TAG_WIDTH-1 downto 0);
      l_discount_cmd_valid         : out std_logic;
      l_discount_cmd_ready         : in  std_logic;
      l_discount_cmd_firstIdx      : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      l_discount_cmd_lastIdx       : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      l_discount_cmd_ctrl          : out std_logic_vector(L_DISCOUNT_BUS_ADDR_WIDTH-1 downto 0);
      l_discount_cmd_tag           : out std_logic_vector(TAG_WIDTH-1 downto 0);
      l_shipdate_cmd_valid         : out std_logic;
      l_shipdate_cmd_ready         : in  std_logic;
      l_shipdate_cmd_firstIdx      : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      l_shipdate_cmd_lastIdx       : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      l_shipdate_cmd_ctrl          : out std_logic_vector(L_SHIPDATE_BUS_ADDR_WIDTH-1 downto 0);
      l_shipdate_cmd_tag           : out std_logic_vector(TAG_WIDTH-1 downto 0)
    );
  end component;

  component Forecast_l is
    generic (
      INDEX_WIDTH                        : integer := 32;
      TAG_WIDTH                          : integer := 1;
      L_QUANTITY_BUS_ADDR_WIDTH          : integer := 64;
      L_QUANTITY_BUS_DATA_WIDTH          : integer := 512;
      L_QUANTITY_BUS_LEN_WIDTH           : integer := 8;
      L_QUANTITY_BUS_BURST_STEP_LEN      : integer := 1;
      L_QUANTITY_BUS_BURST_MAX_LEN       : integer := 16;
      L_EXTENDEDPRICE_BUS_ADDR_WIDTH     : integer := 64;
      L_EXTENDEDPRICE_BUS_DATA_WIDTH     : integer := 512;
      L_EXTENDEDPRICE_BUS_LEN_WIDTH      : integer := 8;
      L_EXTENDEDPRICE_BUS_BURST_STEP_LEN : integer := 1;
      L_EXTENDEDPRICE_BUS_BURST_MAX_LEN  : integer := 16;
      L_DISCOUNT_BUS_ADDR_WIDTH          : integer := 64;
      L_DISCOUNT_BUS_DATA_WIDTH          : integer := 512;
      L_DISCOUNT_BUS_LEN_WIDTH           : integer := 8;
      L_DISCOUNT_BUS_BURST_STEP_LEN      : integer := 1;
      L_DISCOUNT_BUS_BURST_MAX_LEN       : integer := 16;
      L_SHIPDATE_BUS_ADDR_WIDTH          : integer := 64;
      L_SHIPDATE_BUS_DATA_WIDTH          : integer := 512;
      L_SHIPDATE_BUS_LEN_WIDTH           : integer := 8;
      L_SHIPDATE_BUS_BURST_STEP_LEN      : integer := 1;
      L_SHIPDATE_BUS_BURST_MAX_LEN       : integer := 16
    );
    port (
      bcd_clk                        : in  std_logic;
      bcd_reset                      : in  std_logic;
      kcd_clk                        : in  std_logic;
      kcd_reset                      : in  std_logic;
      l_quantity_valid               : out std_logic;
      l_quantity_ready               : in  std_logic;
      l_quantity_dvalid              : out std_logic;
      l_quantity_last                : out std_logic;
      l_quantity                     : out std_logic_vector(63 downto 0);
      l_quantity_bus_rreq_valid      : out std_logic;
      l_quantity_bus_rreq_ready      : in  std_logic;
      l_quantity_bus_rreq_addr       : out std_logic_vector(L_QUANTITY_BUS_ADDR_WIDTH-1 downto 0);
      l_quantity_bus_rreq_len        : out std_logic_vector(L_QUANTITY_BUS_LEN_WIDTH-1 downto 0);
      l_quantity_bus_rdat_valid      : in  std_logic;
      l_quantity_bus_rdat_ready      : out std_logic;
      l_quantity_bus_rdat_data       : in  std_logic_vector(L_QUANTITY_BUS_DATA_WIDTH-1 downto 0);
      l_quantity_bus_rdat_last       : in  std_logic;
      l_quantity_cmd_valid           : in  std_logic;
      l_quantity_cmd_ready           : out std_logic;
      l_quantity_cmd_firstIdx        : in  std_logic_vector(INDEX_WIDTH-1 downto 0);
      l_quantity_cmd_lastIdx         : in  std_logic_vector(INDEX_WIDTH-1 downto 0);
      l_quantity_cmd_ctrl            : in  std_logic_vector(L_QUANTITY_BUS_ADDR_WIDTH-1 downto 0);
      l_quantity_cmd_tag             : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      l_quantity_unl_valid           : out std_logic;
      l_quantity_unl_ready           : in  std_logic;
      l_quantity_unl_tag             : out std_logic_vector(TAG_WIDTH-1 downto 0);
      l_extendedprice_valid          : out std_logic;
      l_extendedprice_ready          : in  std_logic;
      l_extendedprice_dvalid         : out std_logic;
      l_extendedprice_last           : out std_logic;
      l_extendedprice                : out std_logic_vector(63 downto 0);
      l_extendedprice_bus_rreq_valid : out std_logic;
      l_extendedprice_bus_rreq_ready : in  std_logic;
      l_extendedprice_bus_rreq_addr  : out std_logic_vector(L_EXTENDEDPRICE_BUS_ADDR_WIDTH-1 downto 0);
      l_extendedprice_bus_rreq_len   : out std_logic_vector(L_EXTENDEDPRICE_BUS_LEN_WIDTH-1 downto 0);
      l_extendedprice_bus_rdat_valid : in  std_logic;
      l_extendedprice_bus_rdat_ready : out std_logic;
      l_extendedprice_bus_rdat_data  : in  std_logic_vector(L_EXTENDEDPRICE_BUS_DATA_WIDTH-1 downto 0);
      l_extendedprice_bus_rdat_last  : in  std_logic;
      l_extendedprice_cmd_valid      : in  std_logic;
      l_extendedprice_cmd_ready      : out std_logic;
      l_extendedprice_cmd_firstIdx   : in  std_logic_vector(INDEX_WIDTH-1 downto 0);
      l_extendedprice_cmd_lastIdx    : in  std_logic_vector(INDEX_WIDTH-1 downto 0);
      l_extendedprice_cmd_ctrl       : in  std_logic_vector(L_EXTENDEDPRICE_BUS_ADDR_WIDTH-1 downto 0);
      l_extendedprice_cmd_tag        : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      l_extendedprice_unl_valid      : out std_logic;
      l_extendedprice_unl_ready      : in  std_logic;
      l_extendedprice_unl_tag        : out std_logic_vector(TAG_WIDTH-1 downto 0);
      l_discount_valid               : out std_logic;
      l_discount_ready               : in  std_logic;
      l_discount_dvalid              : out std_logic;
      l_discount_last                : out std_logic;
      l_discount                     : out std_logic_vector(63 downto 0);
      l_discount_bus_rreq_valid      : out std_logic;
      l_discount_bus_rreq_ready      : in  std_logic;
      l_discount_bus_rreq_addr       : out std_logic_vector(L_DISCOUNT_BUS_ADDR_WIDTH-1 downto 0);
      l_discount_bus_rreq_len        : out std_logic_vector(L_DISCOUNT_BUS_LEN_WIDTH-1 downto 0);
      l_discount_bus_rdat_valid      : in  std_logic;
      l_discount_bus_rdat_ready      : out std_logic;
      l_discount_bus_rdat_data       : in  std_logic_vector(L_DISCOUNT_BUS_DATA_WIDTH-1 downto 0);
      l_discount_bus_rdat_last       : in  std_logic;
      l_discount_cmd_valid           : in  std_logic;
      l_discount_cmd_ready           : out std_logic;
      l_discount_cmd_firstIdx        : in  std_logic_vector(INDEX_WIDTH-1 downto 0);
      l_discount_cmd_lastIdx         : in  std_logic_vector(INDEX_WIDTH-1 downto 0);
      l_discount_cmd_ctrl            : in  std_logic_vector(L_DISCOUNT_BUS_ADDR_WIDTH-1 downto 0);
      l_discount_cmd_tag             : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      l_discount_unl_valid           : out std_logic;
      l_discount_unl_ready           : in  std_logic;
      l_discount_unl_tag             : out std_logic_vector(TAG_WIDTH-1 downto 0);
      l_shipdate_valid               : out std_logic;
      l_shipdate_ready               : in  std_logic;
      l_shipdate_dvalid              : out std_logic;
      l_shipdate_last                : out std_logic;
      l_shipdate                     : out std_logic_vector(63 downto 0);
      l_shipdate_bus_rreq_valid      : out std_logic;
      l_shipdate_bus_rreq_ready      : in  std_logic;
      l_shipdate_bus_rreq_addr       : out std_logic_vector(L_SHIPDATE_BUS_ADDR_WIDTH-1 downto 0);
      l_shipdate_bus_rreq_len        : out std_logic_vector(L_SHIPDATE_BUS_LEN_WIDTH-1 downto 0);
      l_shipdate_bus_rdat_valid      : in  std_logic;
      l_shipdate_bus_rdat_ready      : out std_logic;
      l_shipdate_bus_rdat_data       : in  std_logic_vector(L_SHIPDATE_BUS_DATA_WIDTH-1 downto 0);
      l_shipdate_bus_rdat_last       : in  std_logic;
      l_shipdate_cmd_valid           : in  std_logic;
      l_shipdate_cmd_ready           : out std_logic;
      l_shipdate_cmd_firstIdx        : in  std_logic_vector(INDEX_WIDTH-1 downto 0);
      l_shipdate_cmd_lastIdx         : in  std_logic_vector(INDEX_WIDTH-1 downto 0);
      l_shipdate_cmd_ctrl            : in  std_logic_vector(L_SHIPDATE_BUS_ADDR_WIDTH-1 downto 0);
      l_shipdate_cmd_tag             : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      l_shipdate_unl_valid           : out std_logic;
      l_shipdate_unl_ready           : in  std_logic;
      l_shipdate_unl_tag             : out std_logic_vector(TAG_WIDTH-1 downto 0)
    );
  end component;

  signal Forecast_Nucleus_inst_mmio_awvalid                 : std_logic;
  signal Forecast_Nucleus_inst_mmio_awready                 : std_logic;
  signal Forecast_Nucleus_inst_mmio_awaddr                  : std_logic_vector(31 downto 0);
  signal Forecast_Nucleus_inst_mmio_wvalid                  : std_logic;
  signal Forecast_Nucleus_inst_mmio_wready                  : std_logic;
  signal Forecast_Nucleus_inst_mmio_wdata                   : std_logic_vector(31 downto 0);
  signal Forecast_Nucleus_inst_mmio_wstrb                   : std_logic_vector(3 downto 0);
  signal Forecast_Nucleus_inst_mmio_bvalid                  : std_logic;
  signal Forecast_Nucleus_inst_mmio_bready                  : std_logic;
  signal Forecast_Nucleus_inst_mmio_bresp                   : std_logic_vector(1 downto 0);
  signal Forecast_Nucleus_inst_mmio_arvalid                 : std_logic;
  signal Forecast_Nucleus_inst_mmio_arready                 : std_logic;
  signal Forecast_Nucleus_inst_mmio_araddr                  : std_logic_vector(31 downto 0);
  signal Forecast_Nucleus_inst_mmio_rvalid                  : std_logic;
  signal Forecast_Nucleus_inst_mmio_rready                  : std_logic;
  signal Forecast_Nucleus_inst_mmio_rdata                   : std_logic_vector(31 downto 0);
  signal Forecast_Nucleus_inst_mmio_rresp                   : std_logic_vector(1 downto 0);

  signal Forecast_Nucleus_inst_l_quantity_valid             : std_logic;
  signal Forecast_Nucleus_inst_l_quantity_ready             : std_logic;
  signal Forecast_Nucleus_inst_l_quantity_dvalid            : std_logic;
  signal Forecast_Nucleus_inst_l_quantity_last              : std_logic;
  signal Forecast_Nucleus_inst_l_quantity                   : std_logic_vector(63 downto 0);

  signal Forecast_Nucleus_inst_l_extendedprice_valid        : std_logic;
  signal Forecast_Nucleus_inst_l_extendedprice_ready        : std_logic;
  signal Forecast_Nucleus_inst_l_extendedprice_dvalid       : std_logic;
  signal Forecast_Nucleus_inst_l_extendedprice_last         : std_logic;
  signal Forecast_Nucleus_inst_l_extendedprice              : std_logic_vector(63 downto 0);

  signal Forecast_Nucleus_inst_l_discount_valid             : std_logic;
  signal Forecast_Nucleus_inst_l_discount_ready             : std_logic;
  signal Forecast_Nucleus_inst_l_discount_dvalid            : std_logic;
  signal Forecast_Nucleus_inst_l_discount_last              : std_logic;
  signal Forecast_Nucleus_inst_l_discount                   : std_logic_vector(63 downto 0);

  signal Forecast_Nucleus_inst_l_shipdate_valid             : std_logic;
  signal Forecast_Nucleus_inst_l_shipdate_ready             : std_logic;
  signal Forecast_Nucleus_inst_l_shipdate_dvalid            : std_logic;
  signal Forecast_Nucleus_inst_l_shipdate_last              : std_logic;
  signal Forecast_Nucleus_inst_l_shipdate                   : std_logic_vector(63 downto 0);

  signal Forecast_Nucleus_inst_l_quantity_unl_valid         : std_logic;
  signal Forecast_Nucleus_inst_l_quantity_unl_ready         : std_logic;
  signal Forecast_Nucleus_inst_l_quantity_unl_tag           : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal Forecast_Nucleus_inst_l_extendedprice_unl_valid    : std_logic;
  signal Forecast_Nucleus_inst_l_extendedprice_unl_ready    : std_logic;
  signal Forecast_Nucleus_inst_l_extendedprice_unl_tag      : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal Forecast_Nucleus_inst_l_discount_unl_valid         : std_logic;
  signal Forecast_Nucleus_inst_l_discount_unl_ready         : std_logic;
  signal Forecast_Nucleus_inst_l_discount_unl_tag           : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal Forecast_Nucleus_inst_l_shipdate_unl_valid         : std_logic;
  signal Forecast_Nucleus_inst_l_shipdate_unl_ready         : std_logic;
  signal Forecast_Nucleus_inst_l_shipdate_unl_tag           : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal Forecast_Nucleus_inst_l_quantity_cmd_valid         : std_logic;
  signal Forecast_Nucleus_inst_l_quantity_cmd_ready         : std_logic;
  signal Forecast_Nucleus_inst_l_quantity_cmd_firstIdx      : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal Forecast_Nucleus_inst_l_quantity_cmd_lastIdx       : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal Forecast_Nucleus_inst_l_quantity_cmd_ctrl          : std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
  signal Forecast_Nucleus_inst_l_quantity_cmd_tag           : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal Forecast_Nucleus_inst_l_extendedprice_cmd_valid    : std_logic;
  signal Forecast_Nucleus_inst_l_extendedprice_cmd_ready    : std_logic;
  signal Forecast_Nucleus_inst_l_extendedprice_cmd_firstIdx : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal Forecast_Nucleus_inst_l_extendedprice_cmd_lastIdx  : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal Forecast_Nucleus_inst_l_extendedprice_cmd_ctrl     : std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
  signal Forecast_Nucleus_inst_l_extendedprice_cmd_tag      : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal Forecast_Nucleus_inst_l_discount_cmd_valid         : std_logic;
  signal Forecast_Nucleus_inst_l_discount_cmd_ready         : std_logic;
  signal Forecast_Nucleus_inst_l_discount_cmd_firstIdx      : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal Forecast_Nucleus_inst_l_discount_cmd_lastIdx       : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal Forecast_Nucleus_inst_l_discount_cmd_ctrl          : std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
  signal Forecast_Nucleus_inst_l_discount_cmd_tag           : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal Forecast_Nucleus_inst_l_shipdate_cmd_valid         : std_logic;
  signal Forecast_Nucleus_inst_l_shipdate_cmd_ready         : std_logic;
  signal Forecast_Nucleus_inst_l_shipdate_cmd_firstIdx      : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal Forecast_Nucleus_inst_l_shipdate_cmd_lastIdx       : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal Forecast_Nucleus_inst_l_shipdate_cmd_ctrl          : std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
  signal Forecast_Nucleus_inst_l_shipdate_cmd_tag           : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal Forecast_l_inst_l_quantity_valid                   : std_logic;
  signal Forecast_l_inst_l_quantity_ready                   : std_logic;
  signal Forecast_l_inst_l_quantity_dvalid                  : std_logic;
  signal Forecast_l_inst_l_quantity_last                    : std_logic;
  signal Forecast_l_inst_l_quantity                         : std_logic_vector(63 downto 0);

  signal Forecast_l_inst_l_quantity_bus_rreq_valid          : std_logic;
  signal Forecast_l_inst_l_quantity_bus_rreq_ready          : std_logic;
  signal Forecast_l_inst_l_quantity_bus_rreq_addr           : std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
  signal Forecast_l_inst_l_quantity_bus_rreq_len            : std_logic_vector(BUS_LEN_WIDTH-1 downto 0);
  signal Forecast_l_inst_l_quantity_bus_rdat_valid          : std_logic;
  signal Forecast_l_inst_l_quantity_bus_rdat_ready          : std_logic;
  signal Forecast_l_inst_l_quantity_bus_rdat_data           : std_logic_vector(BUS_DATA_WIDTH-1 downto 0);
  signal Forecast_l_inst_l_quantity_bus_rdat_last           : std_logic;

  signal Forecast_l_inst_l_quantity_cmd_valid               : std_logic;
  signal Forecast_l_inst_l_quantity_cmd_ready               : std_logic;
  signal Forecast_l_inst_l_quantity_cmd_firstIdx            : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal Forecast_l_inst_l_quantity_cmd_lastIdx             : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal Forecast_l_inst_l_quantity_cmd_ctrl                : std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
  signal Forecast_l_inst_l_quantity_cmd_tag                 : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal Forecast_l_inst_l_quantity_unl_valid               : std_logic;
  signal Forecast_l_inst_l_quantity_unl_ready               : std_logic;
  signal Forecast_l_inst_l_quantity_unl_tag                 : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal Forecast_l_inst_l_extendedprice_valid              : std_logic;
  signal Forecast_l_inst_l_extendedprice_ready              : std_logic;
  signal Forecast_l_inst_l_extendedprice_dvalid             : std_logic;
  signal Forecast_l_inst_l_extendedprice_last               : std_logic;
  signal Forecast_l_inst_l_extendedprice                    : std_logic_vector(63 downto 0);

  signal Forecast_l_inst_l_extendedprice_bus_rreq_valid     : std_logic;
  signal Forecast_l_inst_l_extendedprice_bus_rreq_ready     : std_logic;
  signal Forecast_l_inst_l_extendedprice_bus_rreq_addr      : std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
  signal Forecast_l_inst_l_extendedprice_bus_rreq_len       : std_logic_vector(BUS_LEN_WIDTH-1 downto 0);
  signal Forecast_l_inst_l_extendedprice_bus_rdat_valid     : std_logic;
  signal Forecast_l_inst_l_extendedprice_bus_rdat_ready     : std_logic;
  signal Forecast_l_inst_l_extendedprice_bus_rdat_data      : std_logic_vector(BUS_DATA_WIDTH-1 downto 0);
  signal Forecast_l_inst_l_extendedprice_bus_rdat_last      : std_logic;

  signal Forecast_l_inst_l_extendedprice_cmd_valid          : std_logic;
  signal Forecast_l_inst_l_extendedprice_cmd_ready          : std_logic;
  signal Forecast_l_inst_l_extendedprice_cmd_firstIdx       : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal Forecast_l_inst_l_extendedprice_cmd_lastIdx        : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal Forecast_l_inst_l_extendedprice_cmd_ctrl           : std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
  signal Forecast_l_inst_l_extendedprice_cmd_tag            : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal Forecast_l_inst_l_extendedprice_unl_valid          : std_logic;
  signal Forecast_l_inst_l_extendedprice_unl_ready          : std_logic;
  signal Forecast_l_inst_l_extendedprice_unl_tag            : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal Forecast_l_inst_l_discount_valid                   : std_logic;
  signal Forecast_l_inst_l_discount_ready                   : std_logic;
  signal Forecast_l_inst_l_discount_dvalid                  : std_logic;
  signal Forecast_l_inst_l_discount_last                    : std_logic;
  signal Forecast_l_inst_l_discount                         : std_logic_vector(63 downto 0);

  signal Forecast_l_inst_l_discount_bus_rreq_valid          : std_logic;
  signal Forecast_l_inst_l_discount_bus_rreq_ready          : std_logic;
  signal Forecast_l_inst_l_discount_bus_rreq_addr           : std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
  signal Forecast_l_inst_l_discount_bus_rreq_len            : std_logic_vector(BUS_LEN_WIDTH-1 downto 0);
  signal Forecast_l_inst_l_discount_bus_rdat_valid          : std_logic;
  signal Forecast_l_inst_l_discount_bus_rdat_ready          : std_logic;
  signal Forecast_l_inst_l_discount_bus_rdat_data           : std_logic_vector(BUS_DATA_WIDTH-1 downto 0);
  signal Forecast_l_inst_l_discount_bus_rdat_last           : std_logic;

  signal Forecast_l_inst_l_discount_cmd_valid               : std_logic;
  signal Forecast_l_inst_l_discount_cmd_ready               : std_logic;
  signal Forecast_l_inst_l_discount_cmd_firstIdx            : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal Forecast_l_inst_l_discount_cmd_lastIdx             : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal Forecast_l_inst_l_discount_cmd_ctrl                : std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
  signal Forecast_l_inst_l_discount_cmd_tag                 : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal Forecast_l_inst_l_discount_unl_valid               : std_logic;
  signal Forecast_l_inst_l_discount_unl_ready               : std_logic;
  signal Forecast_l_inst_l_discount_unl_tag                 : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal Forecast_l_inst_l_shipdate_valid                   : std_logic;
  signal Forecast_l_inst_l_shipdate_ready                   : std_logic;
  signal Forecast_l_inst_l_shipdate_dvalid                  : std_logic;
  signal Forecast_l_inst_l_shipdate_last                    : std_logic;
  signal Forecast_l_inst_l_shipdate                         : std_logic_vector(63 downto 0);

  signal Forecast_l_inst_l_shipdate_bus_rreq_valid          : std_logic;
  signal Forecast_l_inst_l_shipdate_bus_rreq_ready          : std_logic;
  signal Forecast_l_inst_l_shipdate_bus_rreq_addr           : std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
  signal Forecast_l_inst_l_shipdate_bus_rreq_len            : std_logic_vector(BUS_LEN_WIDTH-1 downto 0);
  signal Forecast_l_inst_l_shipdate_bus_rdat_valid          : std_logic;
  signal Forecast_l_inst_l_shipdate_bus_rdat_ready          : std_logic;
  signal Forecast_l_inst_l_shipdate_bus_rdat_data           : std_logic_vector(BUS_DATA_WIDTH-1 downto 0);
  signal Forecast_l_inst_l_shipdate_bus_rdat_last           : std_logic;

  signal Forecast_l_inst_l_shipdate_cmd_valid               : std_logic;
  signal Forecast_l_inst_l_shipdate_cmd_ready               : std_logic;
  signal Forecast_l_inst_l_shipdate_cmd_firstIdx            : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal Forecast_l_inst_l_shipdate_cmd_lastIdx             : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal Forecast_l_inst_l_shipdate_cmd_ctrl                : std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
  signal Forecast_l_inst_l_shipdate_cmd_tag                 : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal Forecast_l_inst_l_shipdate_unl_valid               : std_logic;
  signal Forecast_l_inst_l_shipdate_unl_ready               : std_logic;
  signal Forecast_l_inst_l_shipdate_unl_tag                 : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal RDAW64DW512LW8BS1BM16_inst_mst_rreq_valid          : std_logic;
  signal RDAW64DW512LW8BS1BM16_inst_mst_rreq_ready          : std_logic;
  signal RDAW64DW512LW8BS1BM16_inst_mst_rreq_addr           : std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
  signal RDAW64DW512LW8BS1BM16_inst_mst_rreq_len            : std_logic_vector(BUS_LEN_WIDTH-1 downto 0);
  signal RDAW64DW512LW8BS1BM16_inst_mst_rdat_valid          : std_logic;
  signal RDAW64DW512LW8BS1BM16_inst_mst_rdat_ready          : std_logic;
  signal RDAW64DW512LW8BS1BM16_inst_mst_rdat_data           : std_logic_vector(BUS_DATA_WIDTH-1 downto 0);
  signal RDAW64DW512LW8BS1BM16_inst_mst_rdat_last           : std_logic;

  signal RDAW64DW512LW8BS1BM16_inst_bsv_rreq_valid : std_logic_vector(3 downto 0);
  signal RDAW64DW512LW8BS1BM16_inst_bsv_rreq_ready : std_logic_vector(3 downto 0);
  signal RDAW64DW512LW8BS1BM16_inst_bsv_rreq_addr  : std_logic_vector(4*BUS_ADDR_WIDTH-1 downto 0);
  signal RDAW64DW512LW8BS1BM16_inst_bsv_rreq_len   : std_logic_vector(4*BUS_LEN_WIDTH-1 downto 0);
  signal RDAW64DW512LW8BS1BM16_inst_bsv_rdat_valid : std_logic_vector(3 downto 0);
  signal RDAW64DW512LW8BS1BM16_inst_bsv_rdat_ready : std_logic_vector(3 downto 0);
  signal RDAW64DW512LW8BS1BM16_inst_bsv_rdat_data  : std_logic_vector(4*BUS_DATA_WIDTH-1 downto 0);
  signal RDAW64DW512LW8BS1BM16_inst_bsv_rdat_last  : std_logic_vector(3 downto 0);

begin
  Forecast_Nucleus_inst : Forecast_Nucleus
    generic map (
      INDEX_WIDTH                    => INDEX_WIDTH,
      TAG_WIDTH                      => TAG_WIDTH,
      L_QUANTITY_BUS_ADDR_WIDTH      => BUS_ADDR_WIDTH,
      L_EXTENDEDPRICE_BUS_ADDR_WIDTH => BUS_ADDR_WIDTH,
      L_DISCOUNT_BUS_ADDR_WIDTH      => BUS_ADDR_WIDTH,
      L_SHIPDATE_BUS_ADDR_WIDTH      => BUS_ADDR_WIDTH
    )
    port map (
      kcd_clk                      => kcd_clk,
      kcd_reset                    => kcd_reset,
      mmio_awvalid                 => Forecast_Nucleus_inst_mmio_awvalid,
      mmio_awready                 => Forecast_Nucleus_inst_mmio_awready,
      mmio_awaddr                  => Forecast_Nucleus_inst_mmio_awaddr,
      mmio_wvalid                  => Forecast_Nucleus_inst_mmio_wvalid,
      mmio_wready                  => Forecast_Nucleus_inst_mmio_wready,
      mmio_wdata                   => Forecast_Nucleus_inst_mmio_wdata,
      mmio_wstrb                   => Forecast_Nucleus_inst_mmio_wstrb,
      mmio_bvalid                  => Forecast_Nucleus_inst_mmio_bvalid,
      mmio_bready                  => Forecast_Nucleus_inst_mmio_bready,
      mmio_bresp                   => Forecast_Nucleus_inst_mmio_bresp,
      mmio_arvalid                 => Forecast_Nucleus_inst_mmio_arvalid,
      mmio_arready                 => Forecast_Nucleus_inst_mmio_arready,
      mmio_araddr                  => Forecast_Nucleus_inst_mmio_araddr,
      mmio_rvalid                  => Forecast_Nucleus_inst_mmio_rvalid,
      mmio_rready                  => Forecast_Nucleus_inst_mmio_rready,
      mmio_rdata                   => Forecast_Nucleus_inst_mmio_rdata,
      mmio_rresp                   => Forecast_Nucleus_inst_mmio_rresp,
      l_quantity_valid             => Forecast_Nucleus_inst_l_quantity_valid,
      l_quantity_ready             => Forecast_Nucleus_inst_l_quantity_ready,
      l_quantity_dvalid            => Forecast_Nucleus_inst_l_quantity_dvalid,
      l_quantity_last              => Forecast_Nucleus_inst_l_quantity_last,
      l_quantity                   => Forecast_Nucleus_inst_l_quantity,
      l_extendedprice_valid        => Forecast_Nucleus_inst_l_extendedprice_valid,
      l_extendedprice_ready        => Forecast_Nucleus_inst_l_extendedprice_ready,
      l_extendedprice_dvalid       => Forecast_Nucleus_inst_l_extendedprice_dvalid,
      l_extendedprice_last         => Forecast_Nucleus_inst_l_extendedprice_last,
      l_extendedprice              => Forecast_Nucleus_inst_l_extendedprice,
      l_discount_valid             => Forecast_Nucleus_inst_l_discount_valid,
      l_discount_ready             => Forecast_Nucleus_inst_l_discount_ready,
      l_discount_dvalid            => Forecast_Nucleus_inst_l_discount_dvalid,
      l_discount_last              => Forecast_Nucleus_inst_l_discount_last,
      l_discount                   => Forecast_Nucleus_inst_l_discount,
      l_shipdate_valid             => Forecast_Nucleus_inst_l_shipdate_valid,
      l_shipdate_ready             => Forecast_Nucleus_inst_l_shipdate_ready,
      l_shipdate_dvalid            => Forecast_Nucleus_inst_l_shipdate_dvalid,
      l_shipdate_last              => Forecast_Nucleus_inst_l_shipdate_last,
      l_shipdate                   => Forecast_Nucleus_inst_l_shipdate,
      l_quantity_unl_valid         => Forecast_Nucleus_inst_l_quantity_unl_valid,
      l_quantity_unl_ready         => Forecast_Nucleus_inst_l_quantity_unl_ready,
      l_quantity_unl_tag           => Forecast_Nucleus_inst_l_quantity_unl_tag,
      l_extendedprice_unl_valid    => Forecast_Nucleus_inst_l_extendedprice_unl_valid,
      l_extendedprice_unl_ready    => Forecast_Nucleus_inst_l_extendedprice_unl_ready,
      l_extendedprice_unl_tag      => Forecast_Nucleus_inst_l_extendedprice_unl_tag,
      l_discount_unl_valid         => Forecast_Nucleus_inst_l_discount_unl_valid,
      l_discount_unl_ready         => Forecast_Nucleus_inst_l_discount_unl_ready,
      l_discount_unl_tag           => Forecast_Nucleus_inst_l_discount_unl_tag,
      l_shipdate_unl_valid         => Forecast_Nucleus_inst_l_shipdate_unl_valid,
      l_shipdate_unl_ready         => Forecast_Nucleus_inst_l_shipdate_unl_ready,
      l_shipdate_unl_tag           => Forecast_Nucleus_inst_l_shipdate_unl_tag,
      l_quantity_cmd_valid         => Forecast_Nucleus_inst_l_quantity_cmd_valid,
      l_quantity_cmd_ready         => Forecast_Nucleus_inst_l_quantity_cmd_ready,
      l_quantity_cmd_firstIdx      => Forecast_Nucleus_inst_l_quantity_cmd_firstIdx,
      l_quantity_cmd_lastIdx       => Forecast_Nucleus_inst_l_quantity_cmd_lastIdx,
      l_quantity_cmd_ctrl          => Forecast_Nucleus_inst_l_quantity_cmd_ctrl,
      l_quantity_cmd_tag           => Forecast_Nucleus_inst_l_quantity_cmd_tag,
      l_extendedprice_cmd_valid    => Forecast_Nucleus_inst_l_extendedprice_cmd_valid,
      l_extendedprice_cmd_ready    => Forecast_Nucleus_inst_l_extendedprice_cmd_ready,
      l_extendedprice_cmd_firstIdx => Forecast_Nucleus_inst_l_extendedprice_cmd_firstIdx,
      l_extendedprice_cmd_lastIdx  => Forecast_Nucleus_inst_l_extendedprice_cmd_lastIdx,
      l_extendedprice_cmd_ctrl     => Forecast_Nucleus_inst_l_extendedprice_cmd_ctrl,
      l_extendedprice_cmd_tag      => Forecast_Nucleus_inst_l_extendedprice_cmd_tag,
      l_discount_cmd_valid         => Forecast_Nucleus_inst_l_discount_cmd_valid,
      l_discount_cmd_ready         => Forecast_Nucleus_inst_l_discount_cmd_ready,
      l_discount_cmd_firstIdx      => Forecast_Nucleus_inst_l_discount_cmd_firstIdx,
      l_discount_cmd_lastIdx       => Forecast_Nucleus_inst_l_discount_cmd_lastIdx,
      l_discount_cmd_ctrl          => Forecast_Nucleus_inst_l_discount_cmd_ctrl,
      l_discount_cmd_tag           => Forecast_Nucleus_inst_l_discount_cmd_tag,
      l_shipdate_cmd_valid         => Forecast_Nucleus_inst_l_shipdate_cmd_valid,
      l_shipdate_cmd_ready         => Forecast_Nucleus_inst_l_shipdate_cmd_ready,
      l_shipdate_cmd_firstIdx      => Forecast_Nucleus_inst_l_shipdate_cmd_firstIdx,
      l_shipdate_cmd_lastIdx       => Forecast_Nucleus_inst_l_shipdate_cmd_lastIdx,
      l_shipdate_cmd_ctrl          => Forecast_Nucleus_inst_l_shipdate_cmd_ctrl,
      l_shipdate_cmd_tag           => Forecast_Nucleus_inst_l_shipdate_cmd_tag
    );

  Forecast_l_inst : Forecast_l
    generic map (
      INDEX_WIDTH                        => INDEX_WIDTH,
      TAG_WIDTH                          => TAG_WIDTH,
      L_QUANTITY_BUS_ADDR_WIDTH          => BUS_ADDR_WIDTH,
      L_QUANTITY_BUS_DATA_WIDTH          => BUS_DATA_WIDTH,
      L_QUANTITY_BUS_LEN_WIDTH           => BUS_LEN_WIDTH,
      L_QUANTITY_BUS_BURST_STEP_LEN      => BUS_BURST_STEP_LEN,
      L_QUANTITY_BUS_BURST_MAX_LEN       => BUS_BURST_MAX_LEN,
      L_EXTENDEDPRICE_BUS_ADDR_WIDTH     => BUS_ADDR_WIDTH,
      L_EXTENDEDPRICE_BUS_DATA_WIDTH     => BUS_DATA_WIDTH,
      L_EXTENDEDPRICE_BUS_LEN_WIDTH      => BUS_LEN_WIDTH,
      L_EXTENDEDPRICE_BUS_BURST_STEP_LEN => BUS_BURST_STEP_LEN,
      L_EXTENDEDPRICE_BUS_BURST_MAX_LEN  => BUS_BURST_MAX_LEN,
      L_DISCOUNT_BUS_ADDR_WIDTH          => BUS_ADDR_WIDTH,
      L_DISCOUNT_BUS_DATA_WIDTH          => BUS_DATA_WIDTH,
      L_DISCOUNT_BUS_LEN_WIDTH           => BUS_LEN_WIDTH,
      L_DISCOUNT_BUS_BURST_STEP_LEN      => BUS_BURST_STEP_LEN,
      L_DISCOUNT_BUS_BURST_MAX_LEN       => BUS_BURST_MAX_LEN,
      L_SHIPDATE_BUS_ADDR_WIDTH          => BUS_ADDR_WIDTH,
      L_SHIPDATE_BUS_DATA_WIDTH          => BUS_DATA_WIDTH,
      L_SHIPDATE_BUS_LEN_WIDTH           => BUS_LEN_WIDTH,
      L_SHIPDATE_BUS_BURST_STEP_LEN      => BUS_BURST_STEP_LEN,
      L_SHIPDATE_BUS_BURST_MAX_LEN       => BUS_BURST_MAX_LEN
    )
    port map (
      bcd_clk                        => bcd_clk,
      bcd_reset                      => bcd_reset,
      kcd_clk                        => kcd_clk,
      kcd_reset                      => kcd_reset,
      l_quantity_valid               => Forecast_l_inst_l_quantity_valid,
      l_quantity_ready               => Forecast_l_inst_l_quantity_ready,
      l_quantity_dvalid              => Forecast_l_inst_l_quantity_dvalid,
      l_quantity_last                => Forecast_l_inst_l_quantity_last,
      l_quantity                     => Forecast_l_inst_l_quantity,
      l_quantity_bus_rreq_valid      => Forecast_l_inst_l_quantity_bus_rreq_valid,
      l_quantity_bus_rreq_ready      => Forecast_l_inst_l_quantity_bus_rreq_ready,
      l_quantity_bus_rreq_addr       => Forecast_l_inst_l_quantity_bus_rreq_addr,
      l_quantity_bus_rreq_len        => Forecast_l_inst_l_quantity_bus_rreq_len,
      l_quantity_bus_rdat_valid      => Forecast_l_inst_l_quantity_bus_rdat_valid,
      l_quantity_bus_rdat_ready      => Forecast_l_inst_l_quantity_bus_rdat_ready,
      l_quantity_bus_rdat_data       => Forecast_l_inst_l_quantity_bus_rdat_data,
      l_quantity_bus_rdat_last       => Forecast_l_inst_l_quantity_bus_rdat_last,
      l_quantity_cmd_valid           => Forecast_l_inst_l_quantity_cmd_valid,
      l_quantity_cmd_ready           => Forecast_l_inst_l_quantity_cmd_ready,
      l_quantity_cmd_firstIdx        => Forecast_l_inst_l_quantity_cmd_firstIdx,
      l_quantity_cmd_lastIdx         => Forecast_l_inst_l_quantity_cmd_lastIdx,
      l_quantity_cmd_ctrl            => Forecast_l_inst_l_quantity_cmd_ctrl,
      l_quantity_cmd_tag             => Forecast_l_inst_l_quantity_cmd_tag,
      l_quantity_unl_valid           => Forecast_l_inst_l_quantity_unl_valid,
      l_quantity_unl_ready           => Forecast_l_inst_l_quantity_unl_ready,
      l_quantity_unl_tag             => Forecast_l_inst_l_quantity_unl_tag,
      l_extendedprice_valid          => Forecast_l_inst_l_extendedprice_valid,
      l_extendedprice_ready          => Forecast_l_inst_l_extendedprice_ready,
      l_extendedprice_dvalid         => Forecast_l_inst_l_extendedprice_dvalid,
      l_extendedprice_last           => Forecast_l_inst_l_extendedprice_last,
      l_extendedprice                => Forecast_l_inst_l_extendedprice,
      l_extendedprice_bus_rreq_valid => Forecast_l_inst_l_extendedprice_bus_rreq_valid,
      l_extendedprice_bus_rreq_ready => Forecast_l_inst_l_extendedprice_bus_rreq_ready,
      l_extendedprice_bus_rreq_addr  => Forecast_l_inst_l_extendedprice_bus_rreq_addr,
      l_extendedprice_bus_rreq_len   => Forecast_l_inst_l_extendedprice_bus_rreq_len,
      l_extendedprice_bus_rdat_valid => Forecast_l_inst_l_extendedprice_bus_rdat_valid,
      l_extendedprice_bus_rdat_ready => Forecast_l_inst_l_extendedprice_bus_rdat_ready,
      l_extendedprice_bus_rdat_data  => Forecast_l_inst_l_extendedprice_bus_rdat_data,
      l_extendedprice_bus_rdat_last  => Forecast_l_inst_l_extendedprice_bus_rdat_last,
      l_extendedprice_cmd_valid      => Forecast_l_inst_l_extendedprice_cmd_valid,
      l_extendedprice_cmd_ready      => Forecast_l_inst_l_extendedprice_cmd_ready,
      l_extendedprice_cmd_firstIdx   => Forecast_l_inst_l_extendedprice_cmd_firstIdx,
      l_extendedprice_cmd_lastIdx    => Forecast_l_inst_l_extendedprice_cmd_lastIdx,
      l_extendedprice_cmd_ctrl       => Forecast_l_inst_l_extendedprice_cmd_ctrl,
      l_extendedprice_cmd_tag        => Forecast_l_inst_l_extendedprice_cmd_tag,
      l_extendedprice_unl_valid      => Forecast_l_inst_l_extendedprice_unl_valid,
      l_extendedprice_unl_ready      => Forecast_l_inst_l_extendedprice_unl_ready,
      l_extendedprice_unl_tag        => Forecast_l_inst_l_extendedprice_unl_tag,
      l_discount_valid               => Forecast_l_inst_l_discount_valid,
      l_discount_ready               => Forecast_l_inst_l_discount_ready,
      l_discount_dvalid              => Forecast_l_inst_l_discount_dvalid,
      l_discount_last                => Forecast_l_inst_l_discount_last,
      l_discount                     => Forecast_l_inst_l_discount,
      l_discount_bus_rreq_valid      => Forecast_l_inst_l_discount_bus_rreq_valid,
      l_discount_bus_rreq_ready      => Forecast_l_inst_l_discount_bus_rreq_ready,
      l_discount_bus_rreq_addr       => Forecast_l_inst_l_discount_bus_rreq_addr,
      l_discount_bus_rreq_len        => Forecast_l_inst_l_discount_bus_rreq_len,
      l_discount_bus_rdat_valid      => Forecast_l_inst_l_discount_bus_rdat_valid,
      l_discount_bus_rdat_ready      => Forecast_l_inst_l_discount_bus_rdat_ready,
      l_discount_bus_rdat_data       => Forecast_l_inst_l_discount_bus_rdat_data,
      l_discount_bus_rdat_last       => Forecast_l_inst_l_discount_bus_rdat_last,
      l_discount_cmd_valid           => Forecast_l_inst_l_discount_cmd_valid,
      l_discount_cmd_ready           => Forecast_l_inst_l_discount_cmd_ready,
      l_discount_cmd_firstIdx        => Forecast_l_inst_l_discount_cmd_firstIdx,
      l_discount_cmd_lastIdx         => Forecast_l_inst_l_discount_cmd_lastIdx,
      l_discount_cmd_ctrl            => Forecast_l_inst_l_discount_cmd_ctrl,
      l_discount_cmd_tag             => Forecast_l_inst_l_discount_cmd_tag,
      l_discount_unl_valid           => Forecast_l_inst_l_discount_unl_valid,
      l_discount_unl_ready           => Forecast_l_inst_l_discount_unl_ready,
      l_discount_unl_tag             => Forecast_l_inst_l_discount_unl_tag,
      l_shipdate_valid               => Forecast_l_inst_l_shipdate_valid,
      l_shipdate_ready               => Forecast_l_inst_l_shipdate_ready,
      l_shipdate_dvalid              => Forecast_l_inst_l_shipdate_dvalid,
      l_shipdate_last                => Forecast_l_inst_l_shipdate_last,
      l_shipdate                     => Forecast_l_inst_l_shipdate,
      l_shipdate_bus_rreq_valid      => Forecast_l_inst_l_shipdate_bus_rreq_valid,
      l_shipdate_bus_rreq_ready      => Forecast_l_inst_l_shipdate_bus_rreq_ready,
      l_shipdate_bus_rreq_addr       => Forecast_l_inst_l_shipdate_bus_rreq_addr,
      l_shipdate_bus_rreq_len        => Forecast_l_inst_l_shipdate_bus_rreq_len,
      l_shipdate_bus_rdat_valid      => Forecast_l_inst_l_shipdate_bus_rdat_valid,
      l_shipdate_bus_rdat_ready      => Forecast_l_inst_l_shipdate_bus_rdat_ready,
      l_shipdate_bus_rdat_data       => Forecast_l_inst_l_shipdate_bus_rdat_data,
      l_shipdate_bus_rdat_last       => Forecast_l_inst_l_shipdate_bus_rdat_last,
      l_shipdate_cmd_valid           => Forecast_l_inst_l_shipdate_cmd_valid,
      l_shipdate_cmd_ready           => Forecast_l_inst_l_shipdate_cmd_ready,
      l_shipdate_cmd_firstIdx        => Forecast_l_inst_l_shipdate_cmd_firstIdx,
      l_shipdate_cmd_lastIdx         => Forecast_l_inst_l_shipdate_cmd_lastIdx,
      l_shipdate_cmd_ctrl            => Forecast_l_inst_l_shipdate_cmd_ctrl,
      l_shipdate_cmd_tag             => Forecast_l_inst_l_shipdate_cmd_tag,
      l_shipdate_unl_valid           => Forecast_l_inst_l_shipdate_unl_valid,
      l_shipdate_unl_ready           => Forecast_l_inst_l_shipdate_unl_ready,
      l_shipdate_unl_tag             => Forecast_l_inst_l_shipdate_unl_tag
    );

  RDAW64DW512LW8BS1BM16_inst : BusReadArbiterVec
    generic map (
      BUS_ADDR_WIDTH  => BUS_ADDR_WIDTH,
      BUS_DATA_WIDTH  => BUS_DATA_WIDTH,
      BUS_LEN_WIDTH   => BUS_LEN_WIDTH,
      NUM_SLAVE_PORTS => 4,
      ARB_METHOD      => "RR-STICKY",
      MAX_OUTSTANDING => 4,
      RAM_CONFIG      => "",
      SLV_REQ_SLICES  => true,
      MST_REQ_SLICE   => true,
      MST_DAT_SLICE   => true,
      SLV_DAT_SLICES  => true
    )
    port map (
      bcd_clk        => bcd_clk,
      bcd_reset      => bcd_reset,
      mst_rreq_valid => RDAW64DW512LW8BS1BM16_inst_mst_rreq_valid,
      mst_rreq_ready => RDAW64DW512LW8BS1BM16_inst_mst_rreq_ready,
      mst_rreq_addr  => RDAW64DW512LW8BS1BM16_inst_mst_rreq_addr,
      mst_rreq_len   => RDAW64DW512LW8BS1BM16_inst_mst_rreq_len,
      mst_rdat_valid => RDAW64DW512LW8BS1BM16_inst_mst_rdat_valid,
      mst_rdat_ready => RDAW64DW512LW8BS1BM16_inst_mst_rdat_ready,
      mst_rdat_data  => RDAW64DW512LW8BS1BM16_inst_mst_rdat_data,
      mst_rdat_last  => RDAW64DW512LW8BS1BM16_inst_mst_rdat_last,
      bsv_rreq_valid => RDAW64DW512LW8BS1BM16_inst_bsv_rreq_valid,
      bsv_rreq_ready => RDAW64DW512LW8BS1BM16_inst_bsv_rreq_ready,
      bsv_rreq_len   => RDAW64DW512LW8BS1BM16_inst_bsv_rreq_len,
      bsv_rreq_addr  => RDAW64DW512LW8BS1BM16_inst_bsv_rreq_addr,
      bsv_rdat_valid => RDAW64DW512LW8BS1BM16_inst_bsv_rdat_valid,
      bsv_rdat_ready => RDAW64DW512LW8BS1BM16_inst_bsv_rdat_ready,
      bsv_rdat_last  => RDAW64DW512LW8BS1BM16_inst_bsv_rdat_last,
      bsv_rdat_data  => RDAW64DW512LW8BS1BM16_inst_bsv_rdat_data
    );

  rd_mst_rreq_valid                         <= RDAW64DW512LW8BS1BM16_inst_mst_rreq_valid;
  RDAW64DW512LW8BS1BM16_inst_mst_rreq_ready <= rd_mst_rreq_ready;
  rd_mst_rreq_addr                          <= RDAW64DW512LW8BS1BM16_inst_mst_rreq_addr;
  rd_mst_rreq_len                           <= RDAW64DW512LW8BS1BM16_inst_mst_rreq_len;
  RDAW64DW512LW8BS1BM16_inst_mst_rdat_valid <= rd_mst_rdat_valid;
  rd_mst_rdat_ready                         <= RDAW64DW512LW8BS1BM16_inst_mst_rdat_ready;
  RDAW64DW512LW8BS1BM16_inst_mst_rdat_data  <= rd_mst_rdat_data;
  RDAW64DW512LW8BS1BM16_inst_mst_rdat_last  <= rd_mst_rdat_last;

  Forecast_Nucleus_inst_mmio_awvalid              <= mmio_awvalid;
  mmio_awready                                    <= Forecast_Nucleus_inst_mmio_awready;
  Forecast_Nucleus_inst_mmio_awaddr               <= mmio_awaddr;
  Forecast_Nucleus_inst_mmio_wvalid               <= mmio_wvalid;
  mmio_wready                                     <= Forecast_Nucleus_inst_mmio_wready;
  Forecast_Nucleus_inst_mmio_wdata                <= mmio_wdata;
  Forecast_Nucleus_inst_mmio_wstrb                <= mmio_wstrb;
  mmio_bvalid                                     <= Forecast_Nucleus_inst_mmio_bvalid;
  Forecast_Nucleus_inst_mmio_bready               <= mmio_bready;
  mmio_bresp                                      <= Forecast_Nucleus_inst_mmio_bresp;
  Forecast_Nucleus_inst_mmio_arvalid              <= mmio_arvalid;
  mmio_arready                                    <= Forecast_Nucleus_inst_mmio_arready;
  Forecast_Nucleus_inst_mmio_araddr               <= mmio_araddr;
  mmio_rvalid                                     <= Forecast_Nucleus_inst_mmio_rvalid;
  Forecast_Nucleus_inst_mmio_rready               <= mmio_rready;
  mmio_rdata                                      <= Forecast_Nucleus_inst_mmio_rdata;
  mmio_rresp                                      <= Forecast_Nucleus_inst_mmio_rresp;

  Forecast_Nucleus_inst_l_quantity_valid          <= Forecast_l_inst_l_quantity_valid;
  Forecast_l_inst_l_quantity_ready                <= Forecast_Nucleus_inst_l_quantity_ready;
  Forecast_Nucleus_inst_l_quantity_dvalid         <= Forecast_l_inst_l_quantity_dvalid;
  Forecast_Nucleus_inst_l_quantity_last           <= Forecast_l_inst_l_quantity_last;
  Forecast_Nucleus_inst_l_quantity                <= Forecast_l_inst_l_quantity;

  Forecast_Nucleus_inst_l_extendedprice_valid     <= Forecast_l_inst_l_extendedprice_valid;
  Forecast_l_inst_l_extendedprice_ready           <= Forecast_Nucleus_inst_l_extendedprice_ready;
  Forecast_Nucleus_inst_l_extendedprice_dvalid    <= Forecast_l_inst_l_extendedprice_dvalid;
  Forecast_Nucleus_inst_l_extendedprice_last      <= Forecast_l_inst_l_extendedprice_last;
  Forecast_Nucleus_inst_l_extendedprice           <= Forecast_l_inst_l_extendedprice;

  Forecast_Nucleus_inst_l_discount_valid          <= Forecast_l_inst_l_discount_valid;
  Forecast_l_inst_l_discount_ready                <= Forecast_Nucleus_inst_l_discount_ready;
  Forecast_Nucleus_inst_l_discount_dvalid         <= Forecast_l_inst_l_discount_dvalid;
  Forecast_Nucleus_inst_l_discount_last           <= Forecast_l_inst_l_discount_last;
  Forecast_Nucleus_inst_l_discount                <= Forecast_l_inst_l_discount;

  Forecast_Nucleus_inst_l_shipdate_valid          <= Forecast_l_inst_l_shipdate_valid;
  Forecast_l_inst_l_shipdate_ready                <= Forecast_Nucleus_inst_l_shipdate_ready;
  Forecast_Nucleus_inst_l_shipdate_dvalid         <= Forecast_l_inst_l_shipdate_dvalid;
  Forecast_Nucleus_inst_l_shipdate_last           <= Forecast_l_inst_l_shipdate_last;
  Forecast_Nucleus_inst_l_shipdate                <= Forecast_l_inst_l_shipdate;

  Forecast_Nucleus_inst_l_quantity_unl_valid      <= Forecast_l_inst_l_quantity_unl_valid;
  Forecast_l_inst_l_quantity_unl_ready            <= Forecast_Nucleus_inst_l_quantity_unl_ready;
  Forecast_Nucleus_inst_l_quantity_unl_tag        <= Forecast_l_inst_l_quantity_unl_tag;

  Forecast_Nucleus_inst_l_extendedprice_unl_valid <= Forecast_l_inst_l_extendedprice_unl_valid;
  Forecast_l_inst_l_extendedprice_unl_ready       <= Forecast_Nucleus_inst_l_extendedprice_unl_ready;
  Forecast_Nucleus_inst_l_extendedprice_unl_tag   <= Forecast_l_inst_l_extendedprice_unl_tag;

  Forecast_Nucleus_inst_l_discount_unl_valid      <= Forecast_l_inst_l_discount_unl_valid;
  Forecast_l_inst_l_discount_unl_ready            <= Forecast_Nucleus_inst_l_discount_unl_ready;
  Forecast_Nucleus_inst_l_discount_unl_tag        <= Forecast_l_inst_l_discount_unl_tag;

  Forecast_Nucleus_inst_l_shipdate_unl_valid      <= Forecast_l_inst_l_shipdate_unl_valid;
  Forecast_l_inst_l_shipdate_unl_ready            <= Forecast_Nucleus_inst_l_shipdate_unl_ready;
  Forecast_Nucleus_inst_l_shipdate_unl_tag        <= Forecast_l_inst_l_shipdate_unl_tag;

  Forecast_l_inst_l_quantity_cmd_valid            <= Forecast_Nucleus_inst_l_quantity_cmd_valid;
  Forecast_Nucleus_inst_l_quantity_cmd_ready      <= Forecast_l_inst_l_quantity_cmd_ready;
  Forecast_l_inst_l_quantity_cmd_firstIdx         <= Forecast_Nucleus_inst_l_quantity_cmd_firstIdx;
  Forecast_l_inst_l_quantity_cmd_lastIdx          <= Forecast_Nucleus_inst_l_quantity_cmd_lastIdx;
  Forecast_l_inst_l_quantity_cmd_ctrl             <= Forecast_Nucleus_inst_l_quantity_cmd_ctrl;
  Forecast_l_inst_l_quantity_cmd_tag              <= Forecast_Nucleus_inst_l_quantity_cmd_tag;

  Forecast_l_inst_l_extendedprice_cmd_valid       <= Forecast_Nucleus_inst_l_extendedprice_cmd_valid;
  Forecast_Nucleus_inst_l_extendedprice_cmd_ready <= Forecast_l_inst_l_extendedprice_cmd_ready;
  Forecast_l_inst_l_extendedprice_cmd_firstIdx    <= Forecast_Nucleus_inst_l_extendedprice_cmd_firstIdx;
  Forecast_l_inst_l_extendedprice_cmd_lastIdx     <= Forecast_Nucleus_inst_l_extendedprice_cmd_lastIdx;
  Forecast_l_inst_l_extendedprice_cmd_ctrl        <= Forecast_Nucleus_inst_l_extendedprice_cmd_ctrl;
  Forecast_l_inst_l_extendedprice_cmd_tag         <= Forecast_Nucleus_inst_l_extendedprice_cmd_tag;

  Forecast_l_inst_l_discount_cmd_valid            <= Forecast_Nucleus_inst_l_discount_cmd_valid;
  Forecast_Nucleus_inst_l_discount_cmd_ready      <= Forecast_l_inst_l_discount_cmd_ready;
  Forecast_l_inst_l_discount_cmd_firstIdx         <= Forecast_Nucleus_inst_l_discount_cmd_firstIdx;
  Forecast_l_inst_l_discount_cmd_lastIdx          <= Forecast_Nucleus_inst_l_discount_cmd_lastIdx;
  Forecast_l_inst_l_discount_cmd_ctrl             <= Forecast_Nucleus_inst_l_discount_cmd_ctrl;
  Forecast_l_inst_l_discount_cmd_tag              <= Forecast_Nucleus_inst_l_discount_cmd_tag;

  Forecast_l_inst_l_shipdate_cmd_valid            <= Forecast_Nucleus_inst_l_shipdate_cmd_valid;
  Forecast_Nucleus_inst_l_shipdate_cmd_ready      <= Forecast_l_inst_l_shipdate_cmd_ready;
  Forecast_l_inst_l_shipdate_cmd_firstIdx         <= Forecast_Nucleus_inst_l_shipdate_cmd_firstIdx;
  Forecast_l_inst_l_shipdate_cmd_lastIdx          <= Forecast_Nucleus_inst_l_shipdate_cmd_lastIdx;
  Forecast_l_inst_l_shipdate_cmd_ctrl             <= Forecast_Nucleus_inst_l_shipdate_cmd_ctrl;
  Forecast_l_inst_l_shipdate_cmd_tag              <= Forecast_Nucleus_inst_l_shipdate_cmd_tag;

  RDAW64DW512LW8BS1BM16_inst_bsv_rreq_valid(0)                                                        <= Forecast_l_inst_l_quantity_bus_rreq_valid;
  RDAW64DW512LW8BS1BM16_inst_bsv_rreq_valid(1)                                                        <= Forecast_l_inst_l_extendedprice_bus_rreq_valid;
  RDAW64DW512LW8BS1BM16_inst_bsv_rreq_valid(2)                                                        <= Forecast_l_inst_l_discount_bus_rreq_valid;
  RDAW64DW512LW8BS1BM16_inst_bsv_rreq_valid(3)                                                        <= Forecast_l_inst_l_shipdate_bus_rreq_valid;
  RDAW64DW512LW8BS1BM16_inst_bsv_rreq_len(BUS_LEN_WIDTH-1 downto 0)                                   <= Forecast_l_inst_l_quantity_bus_rreq_len;
  RDAW64DW512LW8BS1BM16_inst_bsv_rreq_len(BUS_LEN_WIDTH+BUS_LEN_WIDTH-1 downto BUS_LEN_WIDTH)         <= Forecast_l_inst_l_extendedprice_bus_rreq_len;
  RDAW64DW512LW8BS1BM16_inst_bsv_rreq_len(BUS_LEN_WIDTH*2+BUS_LEN_WIDTH-1 downto BUS_LEN_WIDTH*2)     <= Forecast_l_inst_l_discount_bus_rreq_len;
  RDAW64DW512LW8BS1BM16_inst_bsv_rreq_len(BUS_LEN_WIDTH*3+BUS_LEN_WIDTH-1 downto BUS_LEN_WIDTH*3)     <= Forecast_l_inst_l_shipdate_bus_rreq_len;
  RDAW64DW512LW8BS1BM16_inst_bsv_rreq_addr(BUS_ADDR_WIDTH-1 downto 0)                                 <= Forecast_l_inst_l_quantity_bus_rreq_addr;
  RDAW64DW512LW8BS1BM16_inst_bsv_rreq_addr(BUS_ADDR_WIDTH+BUS_ADDR_WIDTH-1 downto BUS_ADDR_WIDTH)     <= Forecast_l_inst_l_extendedprice_bus_rreq_addr;
  RDAW64DW512LW8BS1BM16_inst_bsv_rreq_addr(BUS_ADDR_WIDTH*2+BUS_ADDR_WIDTH-1 downto BUS_ADDR_WIDTH*2) <= Forecast_l_inst_l_discount_bus_rreq_addr;
  RDAW64DW512LW8BS1BM16_inst_bsv_rreq_addr(BUS_ADDR_WIDTH*3+BUS_ADDR_WIDTH-1 downto BUS_ADDR_WIDTH*3) <= Forecast_l_inst_l_shipdate_bus_rreq_addr;
  RDAW64DW512LW8BS1BM16_inst_bsv_rdat_ready(0)                                                        <= Forecast_l_inst_l_quantity_bus_rdat_ready;
  RDAW64DW512LW8BS1BM16_inst_bsv_rdat_ready(1)                                                        <= Forecast_l_inst_l_extendedprice_bus_rdat_ready;
  RDAW64DW512LW8BS1BM16_inst_bsv_rdat_ready(2)                                                        <= Forecast_l_inst_l_discount_bus_rdat_ready;
  RDAW64DW512LW8BS1BM16_inst_bsv_rdat_ready(3)                                                        <= Forecast_l_inst_l_shipdate_bus_rdat_ready;
  Forecast_l_inst_l_shipdate_bus_rreq_ready                                                           <= RDAW64DW512LW8BS1BM16_inst_bsv_rreq_ready(3);
  Forecast_l_inst_l_shipdate_bus_rdat_valid                                                           <= RDAW64DW512LW8BS1BM16_inst_bsv_rdat_valid(3);
  Forecast_l_inst_l_shipdate_bus_rdat_last                                                            <= RDAW64DW512LW8BS1BM16_inst_bsv_rdat_last(3);
  Forecast_l_inst_l_shipdate_bus_rdat_data                                                            <= RDAW64DW512LW8BS1BM16_inst_bsv_rdat_data(BUS_DATA_WIDTH*3+BUS_DATA_WIDTH-1 downto BUS_DATA_WIDTH*3);
  Forecast_l_inst_l_quantity_bus_rreq_ready                                                           <= RDAW64DW512LW8BS1BM16_inst_bsv_rreq_ready(0);
  Forecast_l_inst_l_quantity_bus_rdat_valid                                                           <= RDAW64DW512LW8BS1BM16_inst_bsv_rdat_valid(0);
  Forecast_l_inst_l_quantity_bus_rdat_last                                                            <= RDAW64DW512LW8BS1BM16_inst_bsv_rdat_last(0);
  Forecast_l_inst_l_quantity_bus_rdat_data                                                            <= RDAW64DW512LW8BS1BM16_inst_bsv_rdat_data(BUS_DATA_WIDTH-1 downto 0);
  Forecast_l_inst_l_extendedprice_bus_rreq_ready                                                      <= RDAW64DW512LW8BS1BM16_inst_bsv_rreq_ready(1);
  Forecast_l_inst_l_extendedprice_bus_rdat_valid                                                      <= RDAW64DW512LW8BS1BM16_inst_bsv_rdat_valid(1);
  Forecast_l_inst_l_extendedprice_bus_rdat_last                                                       <= RDAW64DW512LW8BS1BM16_inst_bsv_rdat_last(1);
  Forecast_l_inst_l_extendedprice_bus_rdat_data                                                       <= RDAW64DW512LW8BS1BM16_inst_bsv_rdat_data(BUS_DATA_WIDTH+BUS_DATA_WIDTH-1 downto BUS_DATA_WIDTH);
  Forecast_l_inst_l_discount_bus_rreq_ready                                                           <= RDAW64DW512LW8BS1BM16_inst_bsv_rreq_ready(2);
  Forecast_l_inst_l_discount_bus_rdat_valid                                                           <= RDAW64DW512LW8BS1BM16_inst_bsv_rdat_valid(2);
  Forecast_l_inst_l_discount_bus_rdat_last                                                            <= RDAW64DW512LW8BS1BM16_inst_bsv_rdat_last(2);
  Forecast_l_inst_l_discount_bus_rdat_data                                                            <= RDAW64DW512LW8BS1BM16_inst_bsv_rdat_data(BUS_DATA_WIDTH*2+BUS_DATA_WIDTH-1 downto BUS_DATA_WIDTH*2);

end architecture;
