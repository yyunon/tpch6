-- Copyright 2018-2019 Delft University of Technology
--
-- Licensed under the Apache License, Version 2.0 (the "License");
-- you may not use this file except in compliance with the License.
-- You may obtain a copy of the License at
--
--     http://www.apache.org/licenses/LICENSE-2.0
--
-- Unless required by applicable law or agreed to in writing, software
-- distributed under the License is distributed on an "AS IS" BASIS,
-- WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
-- See the License for the specific language governing permissions and
-- limitations under the License.
--
-- This file was generated by Fletchgen. Modify this file at your own risk.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.Array_pkg.all;
use work.mmio_pkg.all;

entity Forecast_Nucleus is
  generic (
    INDEX_WIDTH                    : integer := 32;
    TAG_WIDTH                      : integer := 1;
    L_QUANTITY_BUS_ADDR_WIDTH      : integer := 64;
    L_EXTENDEDPRICE_BUS_ADDR_WIDTH : integer := 64;
    L_DISCOUNT_BUS_ADDR_WIDTH      : integer := 64;
    L_SHIPDATE_BUS_ADDR_WIDTH      : integer := 64
  );
  port (
    kcd_clk                      : in  std_logic;
    kcd_reset                    : in  std_logic;
    mmio_awvalid                 : in  std_logic;
    mmio_awready                 : out std_logic;
    mmio_awaddr                  : in  std_logic_vector(31 downto 0);
    mmio_wvalid                  : in  std_logic;
    mmio_wready                  : out std_logic;
    mmio_wdata                   : in  std_logic_vector(31 downto 0);
    mmio_wstrb                   : in  std_logic_vector(3 downto 0);
    mmio_bvalid                  : out std_logic;
    mmio_bready                  : in  std_logic;
    mmio_bresp                   : out std_logic_vector(1 downto 0);
    mmio_arvalid                 : in  std_logic;
    mmio_arready                 : out std_logic;
    mmio_araddr                  : in  std_logic_vector(31 downto 0);
    mmio_rvalid                  : out std_logic;
    mmio_rready                  : in  std_logic;
    mmio_rdata                   : out std_logic_vector(31 downto 0);
    mmio_rresp                   : out std_logic_vector(1 downto 0);
    l_quantity_valid             : in  std_logic;
    l_quantity_ready             : out std_logic;
    l_quantity_dvalid            : in  std_logic;
    l_quantity_last              : in  std_logic;
    l_quantity                   : in  std_logic_vector(511 downto 0);
    l_quantity_count             : in  std_logic_vector(3 downto 0);
    l_extendedprice_valid        : in  std_logic;
    l_extendedprice_ready        : out std_logic;
    l_extendedprice_dvalid       : in  std_logic;
    l_extendedprice_last         : in  std_logic;
    l_extendedprice              : in  std_logic_vector(511 downto 0);
    l_extendedprice_count        : in  std_logic_vector(3 downto 0);
    l_discount_valid             : in  std_logic;
    l_discount_ready             : out std_logic;
    l_discount_dvalid            : in  std_logic;
    l_discount_last              : in  std_logic;
    l_discount                   : in  std_logic_vector(511 downto 0);
    l_discount_count             : in  std_logic_vector(3 downto 0);
    l_shipdate_valid             : in  std_logic;
    l_shipdate_ready             : out std_logic;
    l_shipdate_dvalid            : in  std_logic;
    l_shipdate_last              : in  std_logic;
    l_shipdate                   : in  std_logic_vector(511 downto 0);
    l_shipdate_count             : in  std_logic_vector(3 downto 0);
    l_quantity_unl_valid         : in  std_logic;
    l_quantity_unl_ready         : out std_logic;
    l_quantity_unl_tag           : in  std_logic_vector(TAG_WIDTH-1 downto 0);
    l_extendedprice_unl_valid    : in  std_logic;
    l_extendedprice_unl_ready    : out std_logic;
    l_extendedprice_unl_tag      : in  std_logic_vector(TAG_WIDTH-1 downto 0);
    l_discount_unl_valid         : in  std_logic;
    l_discount_unl_ready         : out std_logic;
    l_discount_unl_tag           : in  std_logic_vector(TAG_WIDTH-1 downto 0);
    l_shipdate_unl_valid         : in  std_logic;
    l_shipdate_unl_ready         : out std_logic;
    l_shipdate_unl_tag           : in  std_logic_vector(TAG_WIDTH-1 downto 0);
    l_quantity_cmd_valid         : out std_logic;
    l_quantity_cmd_ready         : in  std_logic;
    l_quantity_cmd_firstIdx      : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    l_quantity_cmd_lastIdx       : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    l_quantity_cmd_ctrl          : out std_logic_vector(L_QUANTITY_BUS_ADDR_WIDTH-1 downto 0);
    l_quantity_cmd_tag           : out std_logic_vector(TAG_WIDTH-1 downto 0);
    l_extendedprice_cmd_valid    : out std_logic;
    l_extendedprice_cmd_ready    : in  std_logic;
    l_extendedprice_cmd_firstIdx : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    l_extendedprice_cmd_lastIdx  : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    l_extendedprice_cmd_ctrl     : out std_logic_vector(L_EXTENDEDPRICE_BUS_ADDR_WIDTH-1 downto 0);
    l_extendedprice_cmd_tag      : out std_logic_vector(TAG_WIDTH-1 downto 0);
    l_discount_cmd_valid         : out std_logic;
    l_discount_cmd_ready         : in  std_logic;
    l_discount_cmd_firstIdx      : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    l_discount_cmd_lastIdx       : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    l_discount_cmd_ctrl          : out std_logic_vector(L_DISCOUNT_BUS_ADDR_WIDTH-1 downto 0);
    l_discount_cmd_tag           : out std_logic_vector(TAG_WIDTH-1 downto 0);
    l_shipdate_cmd_valid         : out std_logic;
    l_shipdate_cmd_ready         : in  std_logic;
    l_shipdate_cmd_firstIdx      : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    l_shipdate_cmd_lastIdx       : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    l_shipdate_cmd_ctrl          : out std_logic_vector(L_SHIPDATE_BUS_ADDR_WIDTH-1 downto 0);
    l_shipdate_cmd_tag           : out std_logic_vector(TAG_WIDTH-1 downto 0)
  );
end entity;

architecture Implementation of Forecast_Nucleus is
  component Forecast is
    generic (
      INDEX_WIDTH : integer := 32;
      TAG_WIDTH   : integer := 1
    );
    port (
      kcd_clk                      : in  std_logic;
      kcd_reset                    : in  std_logic;
      l_quantity_valid             : in  std_logic;
      l_quantity_ready             : out std_logic;
      l_quantity_dvalid            : in  std_logic;
      l_quantity_last              : in  std_logic;
      l_quantity                   : in  std_logic_vector(511 downto 0);
      l_quantity_count             : in  std_logic_vector(3 downto 0);
      l_extendedprice_valid        : in  std_logic;
      l_extendedprice_ready        : out std_logic;
      l_extendedprice_dvalid       : in  std_logic;
      l_extendedprice_last         : in  std_logic;
      l_extendedprice              : in  std_logic_vector(511 downto 0);
      l_extendedprice_count        : in  std_logic_vector(3 downto 0);
      l_discount_valid             : in  std_logic;
      l_discount_ready             : out std_logic;
      l_discount_dvalid            : in  std_logic;
      l_discount_last              : in  std_logic;
      l_discount                   : in  std_logic_vector(511 downto 0);
      l_discount_count             : in  std_logic_vector(3 downto 0);
      l_shipdate_valid             : in  std_logic;
      l_shipdate_ready             : out std_logic;
      l_shipdate_dvalid            : in  std_logic;
      l_shipdate_last              : in  std_logic;
      l_shipdate                   : in  std_logic_vector(511 downto 0);
      l_shipdate_count             : in  std_logic_vector(3 downto 0);
      l_quantity_unl_valid         : in  std_logic;
      l_quantity_unl_ready         : out std_logic;
      l_quantity_unl_tag           : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      l_extendedprice_unl_valid    : in  std_logic;
      l_extendedprice_unl_ready    : out std_logic;
      l_extendedprice_unl_tag      : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      l_discount_unl_valid         : in  std_logic;
      l_discount_unl_ready         : out std_logic;
      l_discount_unl_tag           : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      l_shipdate_unl_valid         : in  std_logic;
      l_shipdate_unl_ready         : out std_logic;
      l_shipdate_unl_tag           : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      l_quantity_cmd_valid         : out std_logic;
      l_quantity_cmd_ready         : in  std_logic;
      l_quantity_cmd_firstIdx      : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      l_quantity_cmd_lastIdx       : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      l_quantity_cmd_tag           : out std_logic_vector(TAG_WIDTH-1 downto 0);
      l_extendedprice_cmd_valid    : out std_logic;
      l_extendedprice_cmd_ready    : in  std_logic;
      l_extendedprice_cmd_firstIdx : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      l_extendedprice_cmd_lastIdx  : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      l_extendedprice_cmd_tag      : out std_logic_vector(TAG_WIDTH-1 downto 0);
      l_discount_cmd_valid         : out std_logic;
      l_discount_cmd_ready         : in  std_logic;
      l_discount_cmd_firstIdx      : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      l_discount_cmd_lastIdx       : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      l_discount_cmd_tag           : out std_logic_vector(TAG_WIDTH-1 downto 0);
      l_shipdate_cmd_valid         : out std_logic;
      l_shipdate_cmd_ready         : in  std_logic;
      l_shipdate_cmd_firstIdx      : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      l_shipdate_cmd_lastIdx       : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      l_shipdate_cmd_tag           : out std_logic_vector(TAG_WIDTH-1 downto 0);
      start                        : in  std_logic;
      stop                         : in  std_logic;
      reset                        : in  std_logic;
      idle                         : out std_logic;
      busy                         : out std_logic;
      done                         : out std_logic;
      result                       : out std_logic_vector(63 downto 0);
      l_firstidx                   : in  std_logic_vector(31 downto 0);
      l_lastidx                    : in  std_logic_vector(31 downto 0);
      rhigh                        : out std_logic_vector(31 downto 0);
      rlow                         : out std_logic_vector(31 downto 0)
    );
  end component;

  signal Forecast_inst_l_quantity_valid                     : std_logic;
  signal Forecast_inst_l_quantity_ready                     : std_logic;
  signal Forecast_inst_l_quantity_dvalid                    : std_logic;
  signal Forecast_inst_l_quantity_last                      : std_logic;
  signal Forecast_inst_l_quantity                           : std_logic_vector(511 downto 0);
  signal Forecast_inst_l_quantity_count                     : std_logic_vector(3 downto 0);

  signal Forecast_inst_l_extendedprice_valid                : std_logic;
  signal Forecast_inst_l_extendedprice_ready                : std_logic;
  signal Forecast_inst_l_extendedprice_dvalid               : std_logic;
  signal Forecast_inst_l_extendedprice_last                 : std_logic;
  signal Forecast_inst_l_extendedprice                      : std_logic_vector(511 downto 0);
  signal Forecast_inst_l_extendedprice_count                : std_logic_vector(3 downto 0);

  signal Forecast_inst_l_discount_valid                     : std_logic;
  signal Forecast_inst_l_discount_ready                     : std_logic;
  signal Forecast_inst_l_discount_dvalid                    : std_logic;
  signal Forecast_inst_l_discount_last                      : std_logic;
  signal Forecast_inst_l_discount                           : std_logic_vector(511 downto 0);
  signal Forecast_inst_l_discount_count                     : std_logic_vector(3 downto 0);

  signal Forecast_inst_l_shipdate_valid                     : std_logic;
  signal Forecast_inst_l_shipdate_ready                     : std_logic;
  signal Forecast_inst_l_shipdate_dvalid                    : std_logic;
  signal Forecast_inst_l_shipdate_last                      : std_logic;
  signal Forecast_inst_l_shipdate                           : std_logic_vector(511 downto 0);
  signal Forecast_inst_l_shipdate_count                     : std_logic_vector(3 downto 0);

  signal Forecast_inst_l_quantity_unl_valid                 : std_logic;
  signal Forecast_inst_l_quantity_unl_ready                 : std_logic;
  signal Forecast_inst_l_quantity_unl_tag                   : std_logic_vector(0 downto 0);

  signal Forecast_inst_l_extendedprice_unl_valid            : std_logic;
  signal Forecast_inst_l_extendedprice_unl_ready            : std_logic;
  signal Forecast_inst_l_extendedprice_unl_tag              : std_logic_vector(0 downto 0);

  signal Forecast_inst_l_discount_unl_valid                 : std_logic;
  signal Forecast_inst_l_discount_unl_ready                 : std_logic;
  signal Forecast_inst_l_discount_unl_tag                   : std_logic_vector(0 downto 0);

  signal Forecast_inst_l_shipdate_unl_valid                 : std_logic;
  signal Forecast_inst_l_shipdate_unl_ready                 : std_logic;
  signal Forecast_inst_l_shipdate_unl_tag                   : std_logic_vector(0 downto 0);

  signal Forecast_inst_l_quantity_cmd_valid                 : std_logic;
  signal Forecast_inst_l_quantity_cmd_ready                 : std_logic;
  signal Forecast_inst_l_quantity_cmd_firstIdx              : std_logic_vector(31 downto 0);
  signal Forecast_inst_l_quantity_cmd_lastIdx               : std_logic_vector(31 downto 0);
  signal Forecast_inst_l_quantity_cmd_tag                   : std_logic_vector(0 downto 0);

  signal Forecast_inst_l_extendedprice_cmd_valid            : std_logic;
  signal Forecast_inst_l_extendedprice_cmd_ready            : std_logic;
  signal Forecast_inst_l_extendedprice_cmd_firstIdx         : std_logic_vector(31 downto 0);
  signal Forecast_inst_l_extendedprice_cmd_lastIdx          : std_logic_vector(31 downto 0);
  signal Forecast_inst_l_extendedprice_cmd_tag              : std_logic_vector(0 downto 0);

  signal Forecast_inst_l_discount_cmd_valid                 : std_logic;
  signal Forecast_inst_l_discount_cmd_ready                 : std_logic;
  signal Forecast_inst_l_discount_cmd_firstIdx              : std_logic_vector(31 downto 0);
  signal Forecast_inst_l_discount_cmd_lastIdx               : std_logic_vector(31 downto 0);
  signal Forecast_inst_l_discount_cmd_tag                   : std_logic_vector(0 downto 0);

  signal Forecast_inst_l_shipdate_cmd_valid                 : std_logic;
  signal Forecast_inst_l_shipdate_cmd_ready                 : std_logic;
  signal Forecast_inst_l_shipdate_cmd_firstIdx              : std_logic_vector(31 downto 0);
  signal Forecast_inst_l_shipdate_cmd_lastIdx               : std_logic_vector(31 downto 0);
  signal Forecast_inst_l_shipdate_cmd_tag                   : std_logic_vector(0 downto 0);

  signal Forecast_inst_start                                : std_logic;
  signal Forecast_inst_stop                                 : std_logic;
  signal Forecast_inst_reset                                : std_logic;
  signal Forecast_inst_idle                                 : std_logic;
  signal Forecast_inst_busy                                 : std_logic;
  signal Forecast_inst_done                                 : std_logic;
  signal Forecast_inst_result                               : std_logic_vector(63 downto 0);
  signal Forecast_inst_l_firstidx                           : std_logic_vector(31 downto 0);
  signal Forecast_inst_l_lastidx                            : std_logic_vector(31 downto 0);
  signal Forecast_inst_rhigh                                : std_logic_vector(31 downto 0);
  signal Forecast_inst_rlow                                 : std_logic_vector(31 downto 0);
  signal mmio_inst_f_start_data                             : std_logic;
  signal mmio_inst_f_stop_data                              : std_logic;
  signal mmio_inst_f_reset_data                             : std_logic;
  signal mmio_inst_f_idle_write_data                        : std_logic;
  signal mmio_inst_f_busy_write_data                        : std_logic;
  signal mmio_inst_f_done_write_data                        : std_logic;
  signal mmio_inst_f_result_write_data                      : std_logic_vector(63 downto 0);
  signal mmio_inst_f_l_firstidx_data                        : std_logic_vector(31 downto 0);
  signal mmio_inst_f_l_lastidx_data                         : std_logic_vector(31 downto 0);
  signal mmio_inst_f_l_quantity_values_data                 : std_logic_vector(63 downto 0);
  signal mmio_inst_f_l_extendedprice_values_data            : std_logic_vector(63 downto 0);
  signal mmio_inst_f_l_discount_values_data                 : std_logic_vector(63 downto 0);
  signal mmio_inst_f_l_shipdate_values_data                 : std_logic_vector(63 downto 0);
  signal mmio_inst_f_rhigh_write_data                       : std_logic_vector(31 downto 0);
  signal mmio_inst_f_rlow_write_data                        : std_logic_vector(31 downto 0);
  signal mmio_inst_f_Profile_enable_data                    : std_logic;
  signal mmio_inst_f_Profile_clear_data                     : std_logic;
  signal mmio_inst_mmio_awvalid                             : std_logic;
  signal mmio_inst_mmio_awready                             : std_logic;
  signal mmio_inst_mmio_awaddr                              : std_logic_vector(31 downto 0);
  signal mmio_inst_mmio_wvalid                              : std_logic;
  signal mmio_inst_mmio_wready                              : std_logic;
  signal mmio_inst_mmio_wdata                               : std_logic_vector(31 downto 0);
  signal mmio_inst_mmio_wstrb                               : std_logic_vector(3 downto 0);
  signal mmio_inst_mmio_bvalid                              : std_logic;
  signal mmio_inst_mmio_bready                              : std_logic;
  signal mmio_inst_mmio_bresp                               : std_logic_vector(1 downto 0);
  signal mmio_inst_mmio_arvalid                             : std_logic;
  signal mmio_inst_mmio_arready                             : std_logic;
  signal mmio_inst_mmio_araddr                              : std_logic_vector(31 downto 0);
  signal mmio_inst_mmio_rvalid                              : std_logic;
  signal mmio_inst_mmio_rready                              : std_logic;
  signal mmio_inst_mmio_rdata                               : std_logic_vector(31 downto 0);
  signal mmio_inst_mmio_rresp                               : std_logic_vector(1 downto 0);

  signal l_quantity_cmd_accm_inst_kernel_cmd_valid          : std_logic;
  signal l_quantity_cmd_accm_inst_kernel_cmd_ready          : std_logic;
  signal l_quantity_cmd_accm_inst_kernel_cmd_firstIdx       : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal l_quantity_cmd_accm_inst_kernel_cmd_lastIdx        : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal l_quantity_cmd_accm_inst_kernel_cmd_tag            : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal l_quantity_cmd_accm_inst_nucleus_cmd_valid         : std_logic;
  signal l_quantity_cmd_accm_inst_nucleus_cmd_ready         : std_logic;
  signal l_quantity_cmd_accm_inst_nucleus_cmd_firstIdx      : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal l_quantity_cmd_accm_inst_nucleus_cmd_lastIdx       : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal l_quantity_cmd_accm_inst_nucleus_cmd_ctrl          : std_logic_vector(L_QUANTITY_BUS_ADDR_WIDTH-1 downto 0);
  signal l_quantity_cmd_accm_inst_nucleus_cmd_tag           : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal l_extendedprice_cmd_accm_inst_kernel_cmd_valid     : std_logic;
  signal l_extendedprice_cmd_accm_inst_kernel_cmd_ready     : std_logic;
  signal l_extendedprice_cmd_accm_inst_kernel_cmd_firstIdx  : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal l_extendedprice_cmd_accm_inst_kernel_cmd_lastIdx   : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal l_extendedprice_cmd_accm_inst_kernel_cmd_tag       : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal l_extendedprice_cmd_accm_inst_nucleus_cmd_valid    : std_logic;
  signal l_extendedprice_cmd_accm_inst_nucleus_cmd_ready    : std_logic;
  signal l_extendedprice_cmd_accm_inst_nucleus_cmd_firstIdx : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal l_extendedprice_cmd_accm_inst_nucleus_cmd_lastIdx  : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal l_extendedprice_cmd_accm_inst_nucleus_cmd_ctrl     : std_logic_vector(L_EXTENDEDPRICE_BUS_ADDR_WIDTH-1 downto 0);
  signal l_extendedprice_cmd_accm_inst_nucleus_cmd_tag      : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal l_discount_cmd_accm_inst_kernel_cmd_valid          : std_logic;
  signal l_discount_cmd_accm_inst_kernel_cmd_ready          : std_logic;
  signal l_discount_cmd_accm_inst_kernel_cmd_firstIdx       : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal l_discount_cmd_accm_inst_kernel_cmd_lastIdx        : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal l_discount_cmd_accm_inst_kernel_cmd_tag            : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal l_discount_cmd_accm_inst_nucleus_cmd_valid         : std_logic;
  signal l_discount_cmd_accm_inst_nucleus_cmd_ready         : std_logic;
  signal l_discount_cmd_accm_inst_nucleus_cmd_firstIdx      : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal l_discount_cmd_accm_inst_nucleus_cmd_lastIdx       : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal l_discount_cmd_accm_inst_nucleus_cmd_ctrl          : std_logic_vector(L_DISCOUNT_BUS_ADDR_WIDTH-1 downto 0);
  signal l_discount_cmd_accm_inst_nucleus_cmd_tag           : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal l_shipdate_cmd_accm_inst_kernel_cmd_valid          : std_logic;
  signal l_shipdate_cmd_accm_inst_kernel_cmd_ready          : std_logic;
  signal l_shipdate_cmd_accm_inst_kernel_cmd_firstIdx       : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal l_shipdate_cmd_accm_inst_kernel_cmd_lastIdx        : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal l_shipdate_cmd_accm_inst_kernel_cmd_tag            : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal l_shipdate_cmd_accm_inst_nucleus_cmd_valid         : std_logic;
  signal l_shipdate_cmd_accm_inst_nucleus_cmd_ready         : std_logic;
  signal l_shipdate_cmd_accm_inst_nucleus_cmd_firstIdx      : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal l_shipdate_cmd_accm_inst_nucleus_cmd_lastIdx       : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal l_shipdate_cmd_accm_inst_nucleus_cmd_ctrl          : std_logic_vector(L_SHIPDATE_BUS_ADDR_WIDTH-1 downto 0);
  signal l_shipdate_cmd_accm_inst_nucleus_cmd_tag           : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal l_quantity_cmd_accm_inst_ctrl      : std_logic_vector(L_QUANTITY_BUS_ADDR_WIDTH-1 downto 0);
  signal l_extendedprice_cmd_accm_inst_ctrl : std_logic_vector(L_EXTENDEDPRICE_BUS_ADDR_WIDTH-1 downto 0);
  signal l_discount_cmd_accm_inst_ctrl      : std_logic_vector(L_DISCOUNT_BUS_ADDR_WIDTH-1 downto 0);
  signal l_shipdate_cmd_accm_inst_ctrl      : std_logic_vector(L_SHIPDATE_BUS_ADDR_WIDTH-1 downto 0);

begin
  Forecast_inst : Forecast
    generic map (
      INDEX_WIDTH => 32,
      TAG_WIDTH   => 1
    )
    port map (
      kcd_clk                      => kcd_clk,
      kcd_reset                    => kcd_reset,
      l_quantity_valid             => Forecast_inst_l_quantity_valid,
      l_quantity_ready             => Forecast_inst_l_quantity_ready,
      l_quantity_dvalid            => Forecast_inst_l_quantity_dvalid,
      l_quantity_last              => Forecast_inst_l_quantity_last,
      l_quantity                   => Forecast_inst_l_quantity,
      l_quantity_count             => Forecast_inst_l_quantity_count,
      l_extendedprice_valid        => Forecast_inst_l_extendedprice_valid,
      l_extendedprice_ready        => Forecast_inst_l_extendedprice_ready,
      l_extendedprice_dvalid       => Forecast_inst_l_extendedprice_dvalid,
      l_extendedprice_last         => Forecast_inst_l_extendedprice_last,
      l_extendedprice              => Forecast_inst_l_extendedprice,
      l_extendedprice_count        => Forecast_inst_l_extendedprice_count,
      l_discount_valid             => Forecast_inst_l_discount_valid,
      l_discount_ready             => Forecast_inst_l_discount_ready,
      l_discount_dvalid            => Forecast_inst_l_discount_dvalid,
      l_discount_last              => Forecast_inst_l_discount_last,
      l_discount                   => Forecast_inst_l_discount,
      l_discount_count             => Forecast_inst_l_discount_count,
      l_shipdate_valid             => Forecast_inst_l_shipdate_valid,
      l_shipdate_ready             => Forecast_inst_l_shipdate_ready,
      l_shipdate_dvalid            => Forecast_inst_l_shipdate_dvalid,
      l_shipdate_last              => Forecast_inst_l_shipdate_last,
      l_shipdate                   => Forecast_inst_l_shipdate,
      l_shipdate_count             => Forecast_inst_l_shipdate_count,
      l_quantity_unl_valid         => Forecast_inst_l_quantity_unl_valid,
      l_quantity_unl_ready         => Forecast_inst_l_quantity_unl_ready,
      l_quantity_unl_tag           => Forecast_inst_l_quantity_unl_tag,
      l_extendedprice_unl_valid    => Forecast_inst_l_extendedprice_unl_valid,
      l_extendedprice_unl_ready    => Forecast_inst_l_extendedprice_unl_ready,
      l_extendedprice_unl_tag      => Forecast_inst_l_extendedprice_unl_tag,
      l_discount_unl_valid         => Forecast_inst_l_discount_unl_valid,
      l_discount_unl_ready         => Forecast_inst_l_discount_unl_ready,
      l_discount_unl_tag           => Forecast_inst_l_discount_unl_tag,
      l_shipdate_unl_valid         => Forecast_inst_l_shipdate_unl_valid,
      l_shipdate_unl_ready         => Forecast_inst_l_shipdate_unl_ready,
      l_shipdate_unl_tag           => Forecast_inst_l_shipdate_unl_tag,
      l_quantity_cmd_valid         => Forecast_inst_l_quantity_cmd_valid,
      l_quantity_cmd_ready         => Forecast_inst_l_quantity_cmd_ready,
      l_quantity_cmd_firstIdx      => Forecast_inst_l_quantity_cmd_firstIdx,
      l_quantity_cmd_lastIdx       => Forecast_inst_l_quantity_cmd_lastIdx,
      l_quantity_cmd_tag           => Forecast_inst_l_quantity_cmd_tag,
      l_extendedprice_cmd_valid    => Forecast_inst_l_extendedprice_cmd_valid,
      l_extendedprice_cmd_ready    => Forecast_inst_l_extendedprice_cmd_ready,
      l_extendedprice_cmd_firstIdx => Forecast_inst_l_extendedprice_cmd_firstIdx,
      l_extendedprice_cmd_lastIdx  => Forecast_inst_l_extendedprice_cmd_lastIdx,
      l_extendedprice_cmd_tag      => Forecast_inst_l_extendedprice_cmd_tag,
      l_discount_cmd_valid         => Forecast_inst_l_discount_cmd_valid,
      l_discount_cmd_ready         => Forecast_inst_l_discount_cmd_ready,
      l_discount_cmd_firstIdx      => Forecast_inst_l_discount_cmd_firstIdx,
      l_discount_cmd_lastIdx       => Forecast_inst_l_discount_cmd_lastIdx,
      l_discount_cmd_tag           => Forecast_inst_l_discount_cmd_tag,
      l_shipdate_cmd_valid         => Forecast_inst_l_shipdate_cmd_valid,
      l_shipdate_cmd_ready         => Forecast_inst_l_shipdate_cmd_ready,
      l_shipdate_cmd_firstIdx      => Forecast_inst_l_shipdate_cmd_firstIdx,
      l_shipdate_cmd_lastIdx       => Forecast_inst_l_shipdate_cmd_lastIdx,
      l_shipdate_cmd_tag           => Forecast_inst_l_shipdate_cmd_tag,
      start                        => Forecast_inst_start,
      stop                         => Forecast_inst_stop,
      reset                        => Forecast_inst_reset,
      idle                         => Forecast_inst_idle,
      busy                         => Forecast_inst_busy,
      done                         => Forecast_inst_done,
      result                       => Forecast_inst_result,
      l_firstidx                   => Forecast_inst_l_firstidx,
      l_lastidx                    => Forecast_inst_l_lastidx,
      rhigh                        => Forecast_inst_rhigh,
      rlow                         => Forecast_inst_rlow
    );

  mmio_inst : mmio
    port map (
      kcd_clk                       => kcd_clk,
      kcd_reset                     => kcd_reset,
      f_start_data                  => mmio_inst_f_start_data,
      f_stop_data                   => mmio_inst_f_stop_data,
      f_reset_data                  => mmio_inst_f_reset_data,
      f_idle_write_data             => mmio_inst_f_idle_write_data,
      f_busy_write_data             => mmio_inst_f_busy_write_data,
      f_done_write_data             => mmio_inst_f_done_write_data,
      f_result_write_data           => mmio_inst_f_result_write_data,
      f_l_firstidx_data             => mmio_inst_f_l_firstidx_data,
      f_l_lastidx_data              => mmio_inst_f_l_lastidx_data,
      f_l_quantity_values_data      => mmio_inst_f_l_quantity_values_data,
      f_l_extendedprice_values_data => mmio_inst_f_l_extendedprice_values_data,
      f_l_discount_values_data      => mmio_inst_f_l_discount_values_data,
      f_l_shipdate_values_data      => mmio_inst_f_l_shipdate_values_data,
      f_rhigh_write_data            => mmio_inst_f_rhigh_write_data,
      f_rlow_write_data             => mmio_inst_f_rlow_write_data,
      mmio_awvalid                  => mmio_inst_mmio_awvalid,
      mmio_awready                  => mmio_inst_mmio_awready,
      mmio_awaddr                   => mmio_inst_mmio_awaddr,
      mmio_wvalid                   => mmio_inst_mmio_wvalid,
      mmio_wready                   => mmio_inst_mmio_wready,
      mmio_wdata                    => mmio_inst_mmio_wdata,
      mmio_wstrb                    => mmio_inst_mmio_wstrb,
      mmio_bvalid                   => mmio_inst_mmio_bvalid,
      mmio_bready                   => mmio_inst_mmio_bready,
      mmio_bresp                    => mmio_inst_mmio_bresp,
      mmio_arvalid                  => mmio_inst_mmio_arvalid,
      mmio_arready                  => mmio_inst_mmio_arready,
      mmio_araddr                   => mmio_inst_mmio_araddr,
      mmio_rvalid                   => mmio_inst_mmio_rvalid,
      mmio_rready                   => mmio_inst_mmio_rready,
      mmio_rdata                    => mmio_inst_mmio_rdata,
      mmio_rresp                    => mmio_inst_mmio_rresp
    );

  l_quantity_cmd_accm_inst : ArrayCmdCtrlMerger
    generic map (
      NUM_ADDR       => 1,
      BUS_ADDR_WIDTH => L_QUANTITY_BUS_ADDR_WIDTH,
      INDEX_WIDTH    => INDEX_WIDTH,
      TAG_WIDTH      => TAG_WIDTH
    )
    port map (
      kernel_cmd_valid     => l_quantity_cmd_accm_inst_kernel_cmd_valid,
      kernel_cmd_ready     => l_quantity_cmd_accm_inst_kernel_cmd_ready,
      kernel_cmd_firstIdx  => l_quantity_cmd_accm_inst_kernel_cmd_firstIdx,
      kernel_cmd_lastIdx   => l_quantity_cmd_accm_inst_kernel_cmd_lastIdx,
      kernel_cmd_tag       => l_quantity_cmd_accm_inst_kernel_cmd_tag,
      nucleus_cmd_valid    => l_quantity_cmd_accm_inst_nucleus_cmd_valid,
      nucleus_cmd_ready    => l_quantity_cmd_accm_inst_nucleus_cmd_ready,
      nucleus_cmd_firstIdx => l_quantity_cmd_accm_inst_nucleus_cmd_firstIdx,
      nucleus_cmd_lastIdx  => l_quantity_cmd_accm_inst_nucleus_cmd_lastIdx,
      nucleus_cmd_ctrl     => l_quantity_cmd_accm_inst_nucleus_cmd_ctrl,
      nucleus_cmd_tag      => l_quantity_cmd_accm_inst_nucleus_cmd_tag,
      ctrl                 => l_quantity_cmd_accm_inst_ctrl
    );

  l_extendedprice_cmd_accm_inst : ArrayCmdCtrlMerger
    generic map (
      NUM_ADDR       => 1,
      BUS_ADDR_WIDTH => L_EXTENDEDPRICE_BUS_ADDR_WIDTH,
      INDEX_WIDTH    => INDEX_WIDTH,
      TAG_WIDTH      => TAG_WIDTH
    )
    port map (
      kernel_cmd_valid     => l_extendedprice_cmd_accm_inst_kernel_cmd_valid,
      kernel_cmd_ready     => l_extendedprice_cmd_accm_inst_kernel_cmd_ready,
      kernel_cmd_firstIdx  => l_extendedprice_cmd_accm_inst_kernel_cmd_firstIdx,
      kernel_cmd_lastIdx   => l_extendedprice_cmd_accm_inst_kernel_cmd_lastIdx,
      kernel_cmd_tag       => l_extendedprice_cmd_accm_inst_kernel_cmd_tag,
      nucleus_cmd_valid    => l_extendedprice_cmd_accm_inst_nucleus_cmd_valid,
      nucleus_cmd_ready    => l_extendedprice_cmd_accm_inst_nucleus_cmd_ready,
      nucleus_cmd_firstIdx => l_extendedprice_cmd_accm_inst_nucleus_cmd_firstIdx,
      nucleus_cmd_lastIdx  => l_extendedprice_cmd_accm_inst_nucleus_cmd_lastIdx,
      nucleus_cmd_ctrl     => l_extendedprice_cmd_accm_inst_nucleus_cmd_ctrl,
      nucleus_cmd_tag      => l_extendedprice_cmd_accm_inst_nucleus_cmd_tag,
      ctrl                 => l_extendedprice_cmd_accm_inst_ctrl
    );

  l_discount_cmd_accm_inst : ArrayCmdCtrlMerger
    generic map (
      NUM_ADDR       => 1,
      BUS_ADDR_WIDTH => L_DISCOUNT_BUS_ADDR_WIDTH,
      INDEX_WIDTH    => INDEX_WIDTH,
      TAG_WIDTH      => TAG_WIDTH
    )
    port map (
      kernel_cmd_valid     => l_discount_cmd_accm_inst_kernel_cmd_valid,
      kernel_cmd_ready     => l_discount_cmd_accm_inst_kernel_cmd_ready,
      kernel_cmd_firstIdx  => l_discount_cmd_accm_inst_kernel_cmd_firstIdx,
      kernel_cmd_lastIdx   => l_discount_cmd_accm_inst_kernel_cmd_lastIdx,
      kernel_cmd_tag       => l_discount_cmd_accm_inst_kernel_cmd_tag,
      nucleus_cmd_valid    => l_discount_cmd_accm_inst_nucleus_cmd_valid,
      nucleus_cmd_ready    => l_discount_cmd_accm_inst_nucleus_cmd_ready,
      nucleus_cmd_firstIdx => l_discount_cmd_accm_inst_nucleus_cmd_firstIdx,
      nucleus_cmd_lastIdx  => l_discount_cmd_accm_inst_nucleus_cmd_lastIdx,
      nucleus_cmd_ctrl     => l_discount_cmd_accm_inst_nucleus_cmd_ctrl,
      nucleus_cmd_tag      => l_discount_cmd_accm_inst_nucleus_cmd_tag,
      ctrl                 => l_discount_cmd_accm_inst_ctrl
    );

  l_shipdate_cmd_accm_inst : ArrayCmdCtrlMerger
    generic map (
      NUM_ADDR       => 1,
      BUS_ADDR_WIDTH => L_SHIPDATE_BUS_ADDR_WIDTH,
      INDEX_WIDTH    => INDEX_WIDTH,
      TAG_WIDTH      => TAG_WIDTH
    )
    port map (
      kernel_cmd_valid     => l_shipdate_cmd_accm_inst_kernel_cmd_valid,
      kernel_cmd_ready     => l_shipdate_cmd_accm_inst_kernel_cmd_ready,
      kernel_cmd_firstIdx  => l_shipdate_cmd_accm_inst_kernel_cmd_firstIdx,
      kernel_cmd_lastIdx   => l_shipdate_cmd_accm_inst_kernel_cmd_lastIdx,
      kernel_cmd_tag       => l_shipdate_cmd_accm_inst_kernel_cmd_tag,
      nucleus_cmd_valid    => l_shipdate_cmd_accm_inst_nucleus_cmd_valid,
      nucleus_cmd_ready    => l_shipdate_cmd_accm_inst_nucleus_cmd_ready,
      nucleus_cmd_firstIdx => l_shipdate_cmd_accm_inst_nucleus_cmd_firstIdx,
      nucleus_cmd_lastIdx  => l_shipdate_cmd_accm_inst_nucleus_cmd_lastIdx,
      nucleus_cmd_ctrl     => l_shipdate_cmd_accm_inst_nucleus_cmd_ctrl,
      nucleus_cmd_tag      => l_shipdate_cmd_accm_inst_nucleus_cmd_tag,
      ctrl                 => l_shipdate_cmd_accm_inst_ctrl
    );

  l_quantity_cmd_valid                            <= l_quantity_cmd_accm_inst_nucleus_cmd_valid;
  l_quantity_cmd_accm_inst_nucleus_cmd_ready      <= l_quantity_cmd_ready;
  l_quantity_cmd_firstIdx                         <= l_quantity_cmd_accm_inst_nucleus_cmd_firstIdx;
  l_quantity_cmd_lastIdx                          <= l_quantity_cmd_accm_inst_nucleus_cmd_lastIdx;
  l_quantity_cmd_ctrl                             <= l_quantity_cmd_accm_inst_nucleus_cmd_ctrl;
  l_quantity_cmd_tag                              <= l_quantity_cmd_accm_inst_nucleus_cmd_tag;

  l_extendedprice_cmd_valid                       <= l_extendedprice_cmd_accm_inst_nucleus_cmd_valid;
  l_extendedprice_cmd_accm_inst_nucleus_cmd_ready <= l_extendedprice_cmd_ready;
  l_extendedprice_cmd_firstIdx                    <= l_extendedprice_cmd_accm_inst_nucleus_cmd_firstIdx;
  l_extendedprice_cmd_lastIdx                     <= l_extendedprice_cmd_accm_inst_nucleus_cmd_lastIdx;
  l_extendedprice_cmd_ctrl                        <= l_extendedprice_cmd_accm_inst_nucleus_cmd_ctrl;
  l_extendedprice_cmd_tag                         <= l_extendedprice_cmd_accm_inst_nucleus_cmd_tag;

  l_discount_cmd_valid                            <= l_discount_cmd_accm_inst_nucleus_cmd_valid;
  l_discount_cmd_accm_inst_nucleus_cmd_ready      <= l_discount_cmd_ready;
  l_discount_cmd_firstIdx                         <= l_discount_cmd_accm_inst_nucleus_cmd_firstIdx;
  l_discount_cmd_lastIdx                          <= l_discount_cmd_accm_inst_nucleus_cmd_lastIdx;
  l_discount_cmd_ctrl                             <= l_discount_cmd_accm_inst_nucleus_cmd_ctrl;
  l_discount_cmd_tag                              <= l_discount_cmd_accm_inst_nucleus_cmd_tag;

  l_shipdate_cmd_valid                            <= l_shipdate_cmd_accm_inst_nucleus_cmd_valid;
  l_shipdate_cmd_accm_inst_nucleus_cmd_ready      <= l_shipdate_cmd_ready;
  l_shipdate_cmd_firstIdx                         <= l_shipdate_cmd_accm_inst_nucleus_cmd_firstIdx;
  l_shipdate_cmd_lastIdx                          <= l_shipdate_cmd_accm_inst_nucleus_cmd_lastIdx;
  l_shipdate_cmd_ctrl                             <= l_shipdate_cmd_accm_inst_nucleus_cmd_ctrl;
  l_shipdate_cmd_tag                              <= l_shipdate_cmd_accm_inst_nucleus_cmd_tag;

  Forecast_inst_l_quantity_valid                    <= l_quantity_valid;
  l_quantity_ready                                  <= Forecast_inst_l_quantity_ready;
  Forecast_inst_l_quantity_dvalid                   <= l_quantity_dvalid;
  Forecast_inst_l_quantity_last                     <= l_quantity_last;
  Forecast_inst_l_quantity                          <= l_quantity;
  Forecast_inst_l_quantity_count                    <= l_quantity_count;

  Forecast_inst_l_extendedprice_valid               <= l_extendedprice_valid;
  l_extendedprice_ready                             <= Forecast_inst_l_extendedprice_ready;
  Forecast_inst_l_extendedprice_dvalid              <= l_extendedprice_dvalid;
  Forecast_inst_l_extendedprice_last                <= l_extendedprice_last;
  Forecast_inst_l_extendedprice                     <= l_extendedprice;
  Forecast_inst_l_extendedprice_count               <= l_extendedprice_count;

  Forecast_inst_l_discount_valid                    <= l_discount_valid;
  l_discount_ready                                  <= Forecast_inst_l_discount_ready;
  Forecast_inst_l_discount_dvalid                   <= l_discount_dvalid;
  Forecast_inst_l_discount_last                     <= l_discount_last;
  Forecast_inst_l_discount                          <= l_discount;
  Forecast_inst_l_discount_count                    <= l_discount_count;

  Forecast_inst_l_shipdate_valid                    <= l_shipdate_valid;
  l_shipdate_ready                                  <= Forecast_inst_l_shipdate_ready;
  Forecast_inst_l_shipdate_dvalid                   <= l_shipdate_dvalid;
  Forecast_inst_l_shipdate_last                     <= l_shipdate_last;
  Forecast_inst_l_shipdate                          <= l_shipdate;
  Forecast_inst_l_shipdate_count                    <= l_shipdate_count;

  Forecast_inst_l_quantity_unl_valid                <= l_quantity_unl_valid;
  l_quantity_unl_ready                              <= Forecast_inst_l_quantity_unl_ready;
  Forecast_inst_l_quantity_unl_tag                  <= l_quantity_unl_tag;

  Forecast_inst_l_extendedprice_unl_valid           <= l_extendedprice_unl_valid;
  l_extendedprice_unl_ready                         <= Forecast_inst_l_extendedprice_unl_ready;
  Forecast_inst_l_extendedprice_unl_tag             <= l_extendedprice_unl_tag;

  Forecast_inst_l_discount_unl_valid                <= l_discount_unl_valid;
  l_discount_unl_ready                              <= Forecast_inst_l_discount_unl_ready;
  Forecast_inst_l_discount_unl_tag                  <= l_discount_unl_tag;

  Forecast_inst_l_shipdate_unl_valid                <= l_shipdate_unl_valid;
  l_shipdate_unl_ready                              <= Forecast_inst_l_shipdate_unl_ready;
  Forecast_inst_l_shipdate_unl_tag                  <= l_shipdate_unl_tag;

  Forecast_inst_start                               <= mmio_inst_f_start_data;
  Forecast_inst_stop                                <= mmio_inst_f_stop_data;
  Forecast_inst_reset                               <= mmio_inst_f_reset_data;
  Forecast_inst_l_firstidx                          <= mmio_inst_f_l_firstidx_data;
  Forecast_inst_l_lastidx                           <= mmio_inst_f_l_lastidx_data;
  mmio_inst_f_idle_write_data                       <= Forecast_inst_idle;
  mmio_inst_f_busy_write_data                       <= Forecast_inst_busy;
  mmio_inst_f_done_write_data                       <= Forecast_inst_done;
  mmio_inst_f_result_write_data                     <= Forecast_inst_result;
  mmio_inst_f_rhigh_write_data                      <= Forecast_inst_rhigh;
  mmio_inst_f_rlow_write_data                       <= Forecast_inst_rlow;
  mmio_inst_mmio_awvalid                            <= mmio_awvalid;
  mmio_awready                                      <= mmio_inst_mmio_awready;
  mmio_inst_mmio_awaddr                             <= mmio_awaddr;
  mmio_inst_mmio_wvalid                             <= mmio_wvalid;
  mmio_wready                                       <= mmio_inst_mmio_wready;
  mmio_inst_mmio_wdata                              <= mmio_wdata;
  mmio_inst_mmio_wstrb                              <= mmio_wstrb;
  mmio_bvalid                                       <= mmio_inst_mmio_bvalid;
  mmio_inst_mmio_bready                             <= mmio_bready;
  mmio_bresp                                        <= mmio_inst_mmio_bresp;
  mmio_inst_mmio_arvalid                            <= mmio_arvalid;
  mmio_arready                                      <= mmio_inst_mmio_arready;
  mmio_inst_mmio_araddr                             <= mmio_araddr;
  mmio_rvalid                                       <= mmio_inst_mmio_rvalid;
  mmio_inst_mmio_rready                             <= mmio_rready;
  mmio_rdata                                        <= mmio_inst_mmio_rdata;
  mmio_rresp                                        <= mmio_inst_mmio_rresp;

  l_quantity_cmd_accm_inst_kernel_cmd_valid         <= Forecast_inst_l_quantity_cmd_valid;
  Forecast_inst_l_quantity_cmd_ready                <= l_quantity_cmd_accm_inst_kernel_cmd_ready;
  l_quantity_cmd_accm_inst_kernel_cmd_firstIdx      <= Forecast_inst_l_quantity_cmd_firstIdx;
  l_quantity_cmd_accm_inst_kernel_cmd_lastIdx       <= Forecast_inst_l_quantity_cmd_lastIdx;
  l_quantity_cmd_accm_inst_kernel_cmd_tag           <= Forecast_inst_l_quantity_cmd_tag;

  l_extendedprice_cmd_accm_inst_kernel_cmd_valid    <= Forecast_inst_l_extendedprice_cmd_valid;
  Forecast_inst_l_extendedprice_cmd_ready           <= l_extendedprice_cmd_accm_inst_kernel_cmd_ready;
  l_extendedprice_cmd_accm_inst_kernel_cmd_firstIdx <= Forecast_inst_l_extendedprice_cmd_firstIdx;
  l_extendedprice_cmd_accm_inst_kernel_cmd_lastIdx  <= Forecast_inst_l_extendedprice_cmd_lastIdx;
  l_extendedprice_cmd_accm_inst_kernel_cmd_tag      <= Forecast_inst_l_extendedprice_cmd_tag;

  l_discount_cmd_accm_inst_kernel_cmd_valid         <= Forecast_inst_l_discount_cmd_valid;
  Forecast_inst_l_discount_cmd_ready                <= l_discount_cmd_accm_inst_kernel_cmd_ready;
  l_discount_cmd_accm_inst_kernel_cmd_firstIdx      <= Forecast_inst_l_discount_cmd_firstIdx;
  l_discount_cmd_accm_inst_kernel_cmd_lastIdx       <= Forecast_inst_l_discount_cmd_lastIdx;
  l_discount_cmd_accm_inst_kernel_cmd_tag           <= Forecast_inst_l_discount_cmd_tag;

  l_shipdate_cmd_accm_inst_kernel_cmd_valid         <= Forecast_inst_l_shipdate_cmd_valid;
  Forecast_inst_l_shipdate_cmd_ready                <= l_shipdate_cmd_accm_inst_kernel_cmd_ready;
  l_shipdate_cmd_accm_inst_kernel_cmd_firstIdx      <= Forecast_inst_l_shipdate_cmd_firstIdx;
  l_shipdate_cmd_accm_inst_kernel_cmd_lastIdx       <= Forecast_inst_l_shipdate_cmd_lastIdx;
  l_shipdate_cmd_accm_inst_kernel_cmd_tag           <= Forecast_inst_l_shipdate_cmd_tag;

  l_quantity_cmd_accm_inst_ctrl(63 downto 0)      <= mmio_inst_f_l_quantity_values_data;
  l_extendedprice_cmd_accm_inst_ctrl(63 downto 0) <= mmio_inst_f_l_extendedprice_values_data;
  l_discount_cmd_accm_inst_ctrl(63 downto 0)      <= mmio_inst_f_l_discount_values_data;
  l_shipdate_cmd_accm_inst_ctrl(63 downto 0)      <= mmio_inst_f_l_shipdate_values_data;

end architecture;
